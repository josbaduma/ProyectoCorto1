`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:46:40 03/28/2016 
// Design Name: 
// Module Name:    ROM_Star 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_Star(
    input [7:0] addr,
    output reg [199:0] data
    );

always @* begin
	case(addr)
		8'h0: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h1: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h2: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h3: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h4: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h5: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h6: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h7: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h8: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h9: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'ha: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'hb: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'hc: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'hd: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'he: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'hf: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h10: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h11: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h12: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h13: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h14: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h15: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h16: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h17: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h18: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h19: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h1a: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h1b: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h1c: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h1d: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h1e: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h1f: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h20: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h21: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h22: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h23: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h24: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h25: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h26: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h27: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h28: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h29: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h2a: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h2b: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h2c: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h2d: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h2e: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h2f: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h30: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h31: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h32: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h33: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h34: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h35: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h36: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h37: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h38: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h39: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h3a: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h3b: data = 200'b00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
		8'h3c: data = 200'b00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000;
		8'h3d: data = 200'b00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000;
		8'h3e: data = 200'b00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000;
		8'h3f: data = 200'b00000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000;
		8'h40: data = 200'b00000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000;
		8'h41: data = 200'b00000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000;
		8'h42: data = 200'b00000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000;
		8'h43: data = 200'b00000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000;
		8'h44: data = 200'b00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000;
		8'h45: data = 200'b00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000;
		8'h46: data = 200'b00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000;
		8'h47: data = 200'b00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000;
		8'h48: data = 200'b00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
		8'h49: data = 200'b00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000;
		8'h4a: data = 200'b00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000;
		8'h4b: data = 200'b00000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000;
		8'h4c: data = 200'b00000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000;
		8'h4d: data = 200'b00000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000;
		8'h4e: data = 200'b00000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000;
		8'h4f: data = 200'b00000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000;
		8'h50: data = 200'b00000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000;
		8'h51: data = 200'b00000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000;
		8'h52: data = 200'b00000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000;
		8'h53: data = 200'b00000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000;
		8'h54: data = 200'b00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
		8'h55: data = 200'b00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
		8'h56: data = 200'b00000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
		8'h57: data = 200'b00000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
		8'h58: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
		8'h59: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000;
		8'h5a: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000;
		8'h5b: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
		8'h5c: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
		8'h5d: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000;
		8'h5e: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000;
		8'h5f: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000;
		8'h60: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000;
		8'h61: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
		8'h62: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
		8'h63: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
		8'h64: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000;
		8'h65: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
		8'h66: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
		8'h67: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
		8'h68: data = 200'b00000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
		8'h69: data = 200'b00000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
		8'h6a: data = 200'b00000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000;
		8'h6b: data = 200'b00000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
		8'h6c: data = 200'b00000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
		8'h6d: data = 200'b00000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000;
		8'h6e: data = 200'b00000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
		8'h6f: data = 200'b00000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
		8'h70: data = 200'b00000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
		8'h71: data = 200'b00000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111100011111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
		8'h72: data = 200'b00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111110000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
		8'h73: data = 200'b00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
		8'h74: data = 200'b00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000;
		8'h75: data = 200'b00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
		8'h76: data = 200'b00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
		8'h77: data = 200'b00000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
		8'h78: data = 200'b00000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
		8'h79: data = 200'b00000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
		8'h7a: data = 200'b00000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
		8'h7b: data = 200'b00000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000;
		8'h7c: data = 200'b00000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000;
		8'h7d: data = 200'b00000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000;
		8'h7e: data = 200'b00000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000;
		8'h7f: data = 200'b00000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000;
		8'h80: data = 200'b00000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000;
		8'h81: data = 200'b00000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000;
		8'h82: data = 200'b00000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000;
		8'h83: data = 200'b00000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000;
		8'h84: data = 200'b00000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000;
		8'h85: data = 200'b00000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000;
		8'h86: data = 200'b00000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000;
		8'h87: data = 200'b00000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000;
		8'h88: data = 200'b00000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000;
		8'h89: data = 200'b00000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000;
		8'h8a: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h8b: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h8c: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h8d: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h8e: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h8f: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h90: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h91: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h92: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h93: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h94: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h95: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase
end

endmodule
