`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:12:09 05/01/2016 
// Design Name: 
// Module Name:    ROM_CardH 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_CardH(
    input clk,
    input [13:0] addr,
    output reg [8:0] data
    );

always @(posedge clk) begin
	case(addr)
		14'h0: data = 9'o0;
		14'h1: data = 9'o0;
		14'h2: data = 9'o0;
		14'h3: data = 9'o0;
		14'h4: data = 9'o0;
		14'h5: data = 9'o0;
		14'h6: data = 9'o0;
		14'h7: data = 9'o0;
		14'h8: data = 9'o0;
		14'h9: data = 9'o0;
		14'ha: data = 9'o0;
		14'hb: data = 9'o0;
		14'hc: data = 9'o0;
		14'hd: data = 9'o0;
		14'he: data = 9'o0;
		14'hf: data = 9'o0;
		14'h10: data = 9'o0;
		14'h11: data = 9'o0;
		14'h12: data = 9'o0;
		14'h13: data = 9'o0;
		14'h14: data = 9'o0;
		14'h15: data = 9'o0;
		14'h16: data = 9'o0;
		14'h17: data = 9'o0;
		14'h18: data = 9'o0;
		14'h19: data = 9'o0;
		14'h1a: data = 9'o0;
		14'h1b: data = 9'o0;
		14'h1c: data = 9'o0;
		14'h1d: data = 9'o0;
		14'h1e: data = 9'o0;
		14'h1f: data = 9'o0;
		14'h20: data = 9'o0;
		14'h21: data = 9'o0;
		14'h22: data = 9'o0;
		14'h23: data = 9'o0;
		14'h24: data = 9'o0;
		14'h25: data = 9'o0;
		14'h26: data = 9'o0;
		14'h27: data = 9'o0;
		14'h28: data = 9'o0;
		14'h29: data = 9'o0;
		14'h2a: data = 9'o0;
		14'h2b: data = 9'o0;
		14'h2c: data = 9'o0;
		14'h2d: data = 9'o0;
		14'h2e: data = 9'o0;
		14'h2f: data = 9'o0;
		14'h30: data = 9'o0;
		14'h31: data = 9'o0;
		14'h32: data = 9'o0;
		14'h33: data = 9'o0;
		14'h34: data = 9'o0;
		14'h35: data = 9'o0;
		14'h36: data = 9'o0;
		14'h37: data = 9'o0;
		14'h38: data = 9'o0;
		14'h39: data = 9'o0;
		14'h3a: data = 9'o0;
		14'h3b: data = 9'o0;
		14'h3c: data = 9'o0;
		14'h3d: data = 9'o0;
		14'h3e: data = 9'o0;
		14'h3f: data = 9'o0;
		14'h40: data = 9'o0;
		14'h41: data = 9'o0;
		14'h42: data = 9'o0;
		14'h43: data = 9'o0;
		14'h44: data = 9'o0;
		14'h45: data = 9'o0;
		14'h46: data = 9'o0;
		14'h47: data = 9'o0;
		14'h48: data = 9'o0;
		14'h49: data = 9'o0;
		14'h4a: data = 9'o0;
		14'h4b: data = 9'o0;
		14'h4c: data = 9'o0;
		14'h4d: data = 9'o0;
		14'h4e: data = 9'o0;
		14'h4f: data = 9'o0;
		14'h50: data = 9'o0;
		14'h51: data = 9'o0;
		14'h52: data = 9'o0;
		14'h53: data = 9'o0;
		14'h54: data = 9'o0;
		14'h55: data = 9'o0;
		14'h56: data = 9'o0;
		14'h57: data = 9'o0;
		14'h58: data = 9'o0;
		14'h59: data = 9'o0;
		14'h5a: data = 9'o0;
		14'h5b: data = 9'o0;
		14'h5c: data = 9'o0;
		14'h5d: data = 9'o0;
		14'h5e: data = 9'o0;
		14'h5f: data = 9'o0;
		14'h60: data = 9'o0;
		14'h61: data = 9'o0;
		14'h62: data = 9'o0;
		14'h63: data = 9'o0;
		14'h64: data = 9'o0;
		14'h65: data = 9'o0;
		14'h66: data = 9'o0;
		14'h67: data = 9'o0;
		14'h68: data = 9'o0;
		14'h69: data = 9'o0;
		14'h6a: data = 9'o0;
		14'h6b: data = 9'o0;
		14'h6c: data = 9'o0;
		14'h6d: data = 9'o0;
		14'h6e: data = 9'o0;
		14'h6f: data = 9'o0;
		14'h70: data = 9'o0;
		14'h71: data = 9'o0;
		14'h72: data = 9'o0;
		14'h73: data = 9'o0;
		14'h74: data = 9'o0;
		14'h75: data = 9'o0;
		14'h76: data = 9'o0;
		14'h77: data = 9'o0;
		14'h78: data = 9'o0;
		14'h79: data = 9'o0;
		14'h7a: data = 9'o0;
		14'h7b: data = 9'o0;
		14'h7c: data = 9'o0;
		14'h7d: data = 9'o0;
		14'h7e: data = 9'o0;
		14'h7f: data = 9'o0;
		14'h80: data = 9'o0;
		14'h81: data = 9'o0;
		14'h82: data = 9'o0;
		14'h83: data = 9'o0;
		14'h84: data = 9'o0;
		14'h85: data = 9'o0;
		14'h86: data = 9'o0;
		14'h87: data = 9'o0;
		14'h88: data = 9'o0;
		14'h89: data = 9'o0;
		14'h8a: data = 9'o0;
		14'h8b: data = 9'o0;
		14'h8c: data = 9'o0;
		14'h8d: data = 9'o0;
		14'h8e: data = 9'o0;
		14'h8f: data = 9'o0;
		14'h90: data = 9'o0;
		14'h91: data = 9'o0;
		14'h92: data = 9'o0;
		14'h93: data = 9'o0;
		14'h94: data = 9'o0;
		14'h95: data = 9'o0;
		14'h96: data = 9'o0;
		14'h97: data = 9'o0;
		14'h98: data = 9'o0;
		14'h99: data = 9'o0;
		14'h9a: data = 9'o0;
		14'h9b: data = 9'o0;
		14'h9c: data = 9'o0;
		14'h9d: data = 9'o0;
		14'h9e: data = 9'o0;
		14'h9f: data = 9'o0;
		14'ha0: data = 9'o0;
		14'ha1: data = 9'o0;
		14'ha2: data = 9'o0;
		14'ha3: data = 9'o0;
		14'ha4: data = 9'o0;
		14'ha5: data = 9'o0;
		14'ha6: data = 9'o0;
		14'ha7: data = 9'o0;
		14'ha8: data = 9'o0;
		14'ha9: data = 9'o0;
		14'haa: data = 9'o0;
		14'hab: data = 9'o0;
		14'hac: data = 9'o0;
		14'had: data = 9'o0;
		14'hae: data = 9'o0;
		14'haf: data = 9'o0;
		14'hb0: data = 9'o0;
		14'hb1: data = 9'o0;
		14'hb2: data = 9'o0;
		14'hb3: data = 9'o0;
		14'hb4: data = 9'o0;
		14'hb5: data = 9'o0;
		14'hb6: data = 9'o0;
		14'hb7: data = 9'o0;
		14'hb8: data = 9'o0;
		14'hb9: data = 9'o0;
		14'hba: data = 9'o0;
		14'hbb: data = 9'o0;
		14'hbc: data = 9'o0;
		14'hbd: data = 9'o0;
		14'hbe: data = 9'o0;
		14'hbf: data = 9'o0;
		14'hc0: data = 9'o0;
		14'hc1: data = 9'o0;
		14'hc2: data = 9'o0;
		14'hc3: data = 9'o0;
		14'hc4: data = 9'o0;
		14'hc5: data = 9'o0;
		14'hc6: data = 9'o0;
		14'hc7: data = 9'o0;
		14'hc8: data = 9'o0;
		14'hc9: data = 9'o0;
		14'hca: data = 9'o0;
		14'hcb: data = 9'o0;
		14'hcc: data = 9'o0;
		14'hcd: data = 9'o0;
		14'hce: data = 9'o0;
		14'hcf: data = 9'o0;
		14'hd0: data = 9'o0;
		14'hd1: data = 9'o0;
		14'hd2: data = 9'o0;
		14'hd3: data = 9'o0;
		14'hd4: data = 9'o0;
		14'hd5: data = 9'o0;
		14'hd6: data = 9'o0;
		14'hd7: data = 9'o0;
		14'hd8: data = 9'o0;
		14'hd9: data = 9'o0;
		14'hda: data = 9'o0;
		14'hdb: data = 9'o0;
		14'hdc: data = 9'o0;
		14'hdd: data = 9'o0;
		14'hde: data = 9'o0;
		14'hdf: data = 9'o0;
		14'he0: data = 9'o0;
		14'he1: data = 9'o0;
		14'he2: data = 9'o0;
		14'he3: data = 9'o0;
		14'he4: data = 9'o0;
		14'he5: data = 9'o0;
		14'he6: data = 9'o0;
		14'he7: data = 9'o0;
		14'he8: data = 9'o0;
		14'he9: data = 9'o0;
		14'hea: data = 9'o0;
		14'heb: data = 9'o0;
		14'hec: data = 9'o0;
		14'hed: data = 9'o0;
		14'hee: data = 9'o0;
		14'hef: data = 9'o0;
		14'hf0: data = 9'o0;
		14'hf1: data = 9'o0;
		14'hf2: data = 9'o0;
		14'hf3: data = 9'o0;
		14'hf4: data = 9'o0;
		14'hf5: data = 9'o0;
		14'hf6: data = 9'o0;
		14'hf7: data = 9'o0;
		14'hf8: data = 9'o0;
		14'hf9: data = 9'o0;
		14'hfa: data = 9'o0;
		14'hfb: data = 9'o0;
		14'hfc: data = 9'o0;
		14'hfd: data = 9'o0;
		14'hfe: data = 9'o0;
		14'hff: data = 9'o0;
		14'h100: data = 9'o0;
		14'h101: data = 9'o0;
		14'h102: data = 9'o0;
		14'h103: data = 9'o0;
		14'h104: data = 9'o0;
		14'h105: data = 9'o0;
		14'h106: data = 9'o0;
		14'h107: data = 9'o0;
		14'h108: data = 9'o0;
		14'h109: data = 9'o0;
		14'h10a: data = 9'o0;
		14'h10b: data = 9'o0;
		14'h10c: data = 9'o0;
		14'h10d: data = 9'o0;
		14'h10e: data = 9'o0;
		14'h10f: data = 9'o0;
		14'h110: data = 9'o0;
		14'h111: data = 9'o0;
		14'h112: data = 9'o0;
		14'h113: data = 9'o0;
		14'h114: data = 9'o0;
		14'h115: data = 9'o0;
		14'h116: data = 9'o0;
		14'h117: data = 9'o0;
		14'h118: data = 9'o0;
		14'h119: data = 9'o0;
		14'h11a: data = 9'o0;
		14'h11b: data = 9'o0;
		14'h11c: data = 9'o0;
		14'h11d: data = 9'o0;
		14'h11e: data = 9'o0;
		14'h11f: data = 9'o0;
		14'h120: data = 9'o0;
		14'h121: data = 9'o0;
		14'h122: data = 9'o0;
		14'h123: data = 9'o0;
		14'h124: data = 9'o0;
		14'h125: data = 9'o0;
		14'h126: data = 9'o0;
		14'h127: data = 9'o0;
		14'h128: data = 9'o0;
		14'h129: data = 9'o0;
		14'h12a: data = 9'o0;
		14'h12b: data = 9'o0;
		14'h12c: data = 9'o0;
		14'h12d: data = 9'o0;
		14'h12e: data = 9'o0;
		14'h12f: data = 9'o0;
		14'h130: data = 9'o0;
		14'h131: data = 9'o0;
		14'h132: data = 9'o0;
		14'h133: data = 9'o0;
		14'h134: data = 9'o0;
		14'h135: data = 9'o0;
		14'h136: data = 9'o0;
		14'h137: data = 9'o0;
		14'h138: data = 9'o0;
		14'h139: data = 9'o0;
		14'h13a: data = 9'o0;
		14'h13b: data = 9'o0;
		14'h13c: data = 9'o0;
		14'h13d: data = 9'o0;
		14'h13e: data = 9'o0;
		14'h13f: data = 9'o0;
		14'h140: data = 9'o0;
		14'h141: data = 9'o0;
		14'h142: data = 9'o0;
		14'h143: data = 9'o0;
		14'h144: data = 9'o0;
		14'h145: data = 9'o0;
		14'h146: data = 9'o0;
		14'h147: data = 9'o0;
		14'h148: data = 9'o0;
		14'h149: data = 9'o0;
		14'h14a: data = 9'o0;
		14'h14b: data = 9'o0;
		14'h14c: data = 9'o0;
		14'h14d: data = 9'o0;
		14'h14e: data = 9'o0;
		14'h14f: data = 9'o0;
		14'h150: data = 9'o0;
		14'h151: data = 9'o0;
		14'h152: data = 9'o0;
		14'h153: data = 9'o0;
		14'h154: data = 9'o0;
		14'h155: data = 9'o0;
		14'h156: data = 9'o0;
		14'h157: data = 9'o0;
		14'h158: data = 9'o0;
		14'h159: data = 9'o0;
		14'h15a: data = 9'o0;
		14'h15b: data = 9'o0;
		14'h15c: data = 9'o0;
		14'h15d: data = 9'o0;
		14'h15e: data = 9'o0;
		14'h15f: data = 9'o0;
		14'h160: data = 9'o0;
		14'h161: data = 9'o0;
		14'h162: data = 9'o0;
		14'h163: data = 9'o0;
		14'h164: data = 9'o0;
		14'h165: data = 9'o0;
		14'h166: data = 9'o0;
		14'h167: data = 9'o0;
		14'h168: data = 9'o0;
		14'h169: data = 9'o0;
		14'h16a: data = 9'o0;
		14'h16b: data = 9'o0;
		14'h16c: data = 9'o0;
		14'h16d: data = 9'o0;
		14'h16e: data = 9'o0;
		14'h16f: data = 9'o0;
		14'h170: data = 9'o0;
		14'h171: data = 9'o0;
		14'h172: data = 9'o0;
		14'h173: data = 9'o0;
		14'h174: data = 9'o0;
		14'h175: data = 9'o0;
		14'h176: data = 9'o0;
		14'h177: data = 9'o0;
		14'h178: data = 9'o0;
		14'h179: data = 9'o0;
		14'h17a: data = 9'o0;
		14'h17b: data = 9'o0;
		14'h17c: data = 9'o0;
		14'h17d: data = 9'o0;
		14'h17e: data = 9'o0;
		14'h17f: data = 9'o0;
		14'h180: data = 9'o0;
		14'h181: data = 9'o0;
		14'h182: data = 9'o0;
		14'h183: data = 9'o0;
		14'h184: data = 9'o0;
		14'h185: data = 9'o0;
		14'h186: data = 9'o0;
		14'h187: data = 9'o0;
		14'h188: data = 9'o0;
		14'h189: data = 9'o0;
		14'h18a: data = 9'o0;
		14'h18b: data = 9'o0;
		14'h18c: data = 9'o0;
		14'h18d: data = 9'o0;
		14'h18e: data = 9'o0;
		14'h18f: data = 9'o0;
		14'h190: data = 9'o0;
		14'h191: data = 9'o0;
		14'h192: data = 9'o0;
		14'h193: data = 9'o0;
		14'h194: data = 9'o0;
		14'h195: data = 9'o0;
		14'h196: data = 9'o0;
		14'h197: data = 9'o0;
		14'h198: data = 9'o0;
		14'h199: data = 9'o0;
		14'h19a: data = 9'o0;
		14'h19b: data = 9'o0;
		14'h19c: data = 9'o0;
		14'h19d: data = 9'o0;
		14'h19e: data = 9'o0;
		14'h19f: data = 9'o0;
		14'h1a0: data = 9'o0;
		14'h1a1: data = 9'o0;
		14'h1a2: data = 9'o0;
		14'h1a3: data = 9'o0;
		14'h1a4: data = 9'o0;
		14'h1a5: data = 9'o0;
		14'h1a6: data = 9'o0;
		14'h1a7: data = 9'o0;
		14'h1a8: data = 9'o0;
		14'h1a9: data = 9'o0;
		14'h1aa: data = 9'o0;
		14'h1ab: data = 9'o0;
		14'h1ac: data = 9'o0;
		14'h1ad: data = 9'o0;
		14'h1ae: data = 9'o0;
		14'h1af: data = 9'o0;
		14'h1b0: data = 9'o0;
		14'h1b1: data = 9'o0;
		14'h1b2: data = 9'o0;
		14'h1b3: data = 9'o0;
		14'h1b4: data = 9'o0;
		14'h1b5: data = 9'o0;
		14'h1b6: data = 9'o0;
		14'h1b7: data = 9'o0;
		14'h1b8: data = 9'o0;
		14'h1b9: data = 9'o0;
		14'h1ba: data = 9'o0;
		14'h1bb: data = 9'o0;
		14'h1bc: data = 9'o0;
		14'h1bd: data = 9'o0;
		14'h1be: data = 9'o0;
		14'h1bf: data = 9'o0;
		14'h1c0: data = 9'o0;
		14'h1c1: data = 9'o0;
		14'h1c2: data = 9'o0;
		14'h1c3: data = 9'o0;
		14'h1c4: data = 9'o0;
		14'h1c5: data = 9'o0;
		14'h1c6: data = 9'o0;
		14'h1c7: data = 9'o0;
		14'h1c8: data = 9'o0;
		14'h1c9: data = 9'o0;
		14'h1ca: data = 9'o0;
		14'h1cb: data = 9'o0;
		14'h1cc: data = 9'o0;
		14'h1cd: data = 9'o0;
		14'h1ce: data = 9'o0;
		14'h1cf: data = 9'o0;
		14'h1d0: data = 9'o0;
		14'h1d1: data = 9'o0;
		14'h1d2: data = 9'o0;
		14'h1d3: data = 9'o0;
		14'h1d4: data = 9'o0;
		14'h1d5: data = 9'o0;
		14'h1d6: data = 9'o0;
		14'h1d7: data = 9'o0;
		14'h1d8: data = 9'o0;
		14'h1d9: data = 9'o0;
		14'h1da: data = 9'o0;
		14'h1db: data = 9'o0;
		14'h1dc: data = 9'o0;
		14'h1dd: data = 9'o0;
		14'h1de: data = 9'o0;
		14'h1df: data = 9'o0;
		14'h1e0: data = 9'o0;
		14'h1e1: data = 9'o0;
		14'h1e2: data = 9'o0;
		14'h1e3: data = 9'o0;
		14'h1e4: data = 9'o0;
		14'h1e5: data = 9'o0;
		14'h1e6: data = 9'o0;
		14'h1e7: data = 9'o0;
		14'h1e8: data = 9'o0;
		14'h1e9: data = 9'o0;
		14'h1ea: data = 9'o0;
		14'h1eb: data = 9'o0;
		14'h1ec: data = 9'o0;
		14'h1ed: data = 9'o0;
		14'h1ee: data = 9'o0;
		14'h1ef: data = 9'o0;
		14'h1f0: data = 9'o0;
		14'h1f1: data = 9'o0;
		14'h1f2: data = 9'o0;
		14'h1f3: data = 9'o0;
		14'h1f4: data = 9'o0;
		14'h1f5: data = 9'o0;
		14'h1f6: data = 9'o0;
		14'h1f7: data = 9'o0;
		14'h1f8: data = 9'o0;
		14'h1f9: data = 9'o0;
		14'h1fa: data = 9'o0;
		14'h1fb: data = 9'o0;
		14'h1fc: data = 9'o0;
		14'h1fd: data = 9'o0;
		14'h1fe: data = 9'o0;
		14'h1ff: data = 9'o0;
		14'h200: data = 9'o0;
		14'h201: data = 9'o0;
		14'h202: data = 9'o0;
		14'h203: data = 9'o0;
		14'h204: data = 9'o0;
		14'h205: data = 9'o0;
		14'h206: data = 9'o0;
		14'h207: data = 9'o0;
		14'h208: data = 9'o0;
		14'h209: data = 9'o0;
		14'h20a: data = 9'o0;
		14'h20b: data = 9'o0;
		14'h20c: data = 9'o0;
		14'h20d: data = 9'o0;
		14'h20e: data = 9'o0;
		14'h20f: data = 9'o0;
		14'h210: data = 9'o0;
		14'h211: data = 9'o0;
		14'h212: data = 9'o0;
		14'h213: data = 9'o0;
		14'h214: data = 9'o0;
		14'h215: data = 9'o0;
		14'h216: data = 9'o0;
		14'h217: data = 9'o0;
		14'h218: data = 9'o0;
		14'h219: data = 9'o0;
		14'h21a: data = 9'o0;
		14'h21b: data = 9'o0;
		14'h21c: data = 9'o0;
		14'h21d: data = 9'o0;
		14'h21e: data = 9'o0;
		14'h21f: data = 9'o0;
		14'h220: data = 9'o0;
		14'h221: data = 9'o0;
		14'h222: data = 9'o0;
		14'h223: data = 9'o0;
		14'h224: data = 9'o0;
		14'h225: data = 9'o0;
		14'h226: data = 9'o0;
		14'h227: data = 9'o0;
		14'h228: data = 9'o0;
		14'h229: data = 9'o0;
		14'h22a: data = 9'o0;
		14'h22b: data = 9'o0;
		14'h22c: data = 9'o0;
		14'h22d: data = 9'o0;
		14'h22e: data = 9'o0;
		14'h22f: data = 9'o0;
		14'h230: data = 9'o0;
		14'h231: data = 9'o0;
		14'h232: data = 9'o0;
		14'h233: data = 9'o0;
		14'h234: data = 9'o0;
		14'h235: data = 9'o0;
		14'h236: data = 9'o0;
		14'h237: data = 9'o0;
		14'h238: data = 9'o0;
		14'h239: data = 9'o0;
		14'h23a: data = 9'o0;
		14'h23b: data = 9'o0;
		14'h23c: data = 9'o0;
		14'h23d: data = 9'o0;
		14'h23e: data = 9'o0;
		14'h23f: data = 9'o0;
		14'h240: data = 9'o0;
		14'h241: data = 9'o0;
		14'h242: data = 9'o0;
		14'h243: data = 9'o0;
		14'h244: data = 9'o0;
		14'h245: data = 9'o0;
		14'h246: data = 9'o0;
		14'h247: data = 9'o0;
		14'h248: data = 9'o0;
		14'h249: data = 9'o0;
		14'h24a: data = 9'o0;
		14'h24b: data = 9'o0;
		14'h24c: data = 9'o0;
		14'h24d: data = 9'o0;
		14'h24e: data = 9'o0;
		14'h24f: data = 9'o0;
		14'h250: data = 9'o0;
		14'h251: data = 9'o0;
		14'h252: data = 9'o0;
		14'h253: data = 9'o0;
		14'h254: data = 9'o0;
		14'h255: data = 9'o0;
		14'h256: data = 9'o0;
		14'h257: data = 9'o0;
		14'h258: data = 9'o0;
		14'h259: data = 9'o0;
		14'h25a: data = 9'o0;
		14'h25b: data = 9'o0;
		14'h25c: data = 9'o0;
		14'h25d: data = 9'o0;
		14'h25e: data = 9'o0;
		14'h25f: data = 9'o0;
		14'h260: data = 9'o0;
		14'h261: data = 9'o0;
		14'h262: data = 9'o0;
		14'h263: data = 9'o0;
		14'h264: data = 9'o0;
		14'h265: data = 9'o0;
		14'h266: data = 9'o0;
		14'h267: data = 9'o0;
		14'h268: data = 9'o0;
		14'h269: data = 9'o0;
		14'h26a: data = 9'o0;
		14'h26b: data = 9'o0;
		14'h26c: data = 9'o0;
		14'h26d: data = 9'o0;
		14'h26e: data = 9'o0;
		14'h26f: data = 9'o0;
		14'h270: data = 9'o0;
		14'h271: data = 9'o0;
		14'h272: data = 9'o0;
		14'h273: data = 9'o0;
		14'h274: data = 9'o0;
		14'h275: data = 9'o0;
		14'h276: data = 9'o0;
		14'h277: data = 9'o0;
		14'h278: data = 9'o0;
		14'h279: data = 9'o0;
		14'h27a: data = 9'o0;
		14'h27b: data = 9'o0;
		14'h27c: data = 9'o0;
		14'h27d: data = 9'o0;
		14'h27e: data = 9'o0;
		14'h27f: data = 9'o0;
		14'h280: data = 9'o0;
		14'h281: data = 9'o0;
		14'h282: data = 9'o0;
		14'h283: data = 9'o0;
		14'h284: data = 9'o0;
		14'h285: data = 9'o0;
		14'h286: data = 9'o0;
		14'h287: data = 9'o0;
		14'h288: data = 9'o0;
		14'h289: data = 9'o0;
		14'h28a: data = 9'o0;
		14'h28b: data = 9'o0;
		14'h28c: data = 9'o0;
		14'h28d: data = 9'o0;
		14'h28e: data = 9'o0;
		14'h28f: data = 9'o0;
		14'h290: data = 9'o0;
		14'h291: data = 9'o0;
		14'h292: data = 9'o0;
		14'h293: data = 9'o0;
		14'h294: data = 9'o0;
		14'h295: data = 9'o0;
		14'h296: data = 9'o0;
		14'h297: data = 9'o0;
		14'h298: data = 9'o0;
		14'h299: data = 9'o0;
		14'h29a: data = 9'o0;
		14'h29b: data = 9'o0;
		14'h29c: data = 9'o0;
		14'h29d: data = 9'o0;
		14'h29e: data = 9'o0;
		14'h29f: data = 9'o0;
		14'h2a0: data = 9'o0;
		14'h2a1: data = 9'o0;
		14'h2a2: data = 9'o0;
		14'h2a3: data = 9'o0;
		14'h2a4: data = 9'o0;
		14'h2a5: data = 9'o0;
		14'h2a6: data = 9'o0;
		14'h2a7: data = 9'o0;
		14'h2a8: data = 9'o0;
		14'h2a9: data = 9'o0;
		14'h2aa: data = 9'o0;
		14'h2ab: data = 9'o0;
		14'h2ac: data = 9'o0;
		14'h2ad: data = 9'o0;
		14'h2ae: data = 9'o0;
		14'h2af: data = 9'o0;
		14'h2b0: data = 9'o0;
		14'h2b1: data = 9'o0;
		14'h2b2: data = 9'o0;
		14'h2b3: data = 9'o0;
		14'h2b4: data = 9'o0;
		14'h2b5: data = 9'o0;
		14'h2b6: data = 9'o0;
		14'h2b7: data = 9'o0;
		14'h2b8: data = 9'o0;
		14'h2b9: data = 9'o0;
		14'h2ba: data = 9'o0;
		14'h2bb: data = 9'o0;
		14'h2bc: data = 9'o0;
		14'h2bd: data = 9'o0;
		14'h2be: data = 9'o0;
		14'h2bf: data = 9'o0;
		14'h2c0: data = 9'o0;
		14'h2c1: data = 9'o0;
		14'h2c2: data = 9'o0;
		14'h2c3: data = 9'o551;
		14'h2c4: data = 9'o652;
		14'h2c5: data = 9'o652;
		14'h2c6: data = 9'o652;
		14'h2c7: data = 9'o652;
		14'h2c8: data = 9'o552;
		14'h2c9: data = 9'o652;
		14'h2ca: data = 9'o652;
		14'h2cb: data = 9'o652;
		14'h2cc: data = 9'o652;
		14'h2cd: data = 9'o551;
		14'h2ce: data = 9'o652;
		14'h2cf: data = 9'o552;
		14'h2d0: data = 9'o652;
		14'h2d1: data = 9'o552;
		14'h2d2: data = 9'o652;
		14'h2d3: data = 9'o652;
		14'h2d4: data = 9'o652;
		14'h2d5: data = 9'o652;
		14'h2d6: data = 9'o552;
		14'h2d7: data = 9'o552;
		14'h2d8: data = 9'o552;
		14'h2d9: data = 9'o552;
		14'h2da: data = 9'o551;
		14'h2db: data = 9'o651;
		14'h2dc: data = 9'o651;
		14'h2dd: data = 9'o651;
		14'h2de: data = 9'o651;
		14'h2df: data = 9'o551;
		14'h2e0: data = 9'o551;
		14'h2e1: data = 9'o551;
		14'h2e2: data = 9'o551;
		14'h2e3: data = 9'o651;
		14'h2e4: data = 9'o651;
		14'h2e5: data = 9'o651;
		14'h2e6: data = 9'o651;
		14'h2e7: data = 9'o551;
		14'h2e8: data = 9'o552;
		14'h2e9: data = 9'o552;
		14'h2ea: data = 9'o552;
		14'h2eb: data = 9'o652;
		14'h2ec: data = 9'o652;
		14'h2ed: data = 9'o652;
		14'h2ee: data = 9'o652;
		14'h2ef: data = 9'o652;
		14'h2f0: data = 9'o652;
		14'h2f1: data = 9'o652;
		14'h2f2: data = 9'o651;
		14'h2f3: data = 9'o652;
		14'h2f4: data = 9'o652;
		14'h2f5: data = 9'o652;
		14'h2f6: data = 9'o552;
		14'h2f7: data = 9'o552;
		14'h2f8: data = 9'o652;
		14'h2f9: data = 9'o652;
		14'h2fa: data = 9'o652;
		14'h2fb: data = 9'o652;
		14'h2fc: data = 9'o552;
		14'h2fd: data = 9'o652;
		14'h2fe: data = 9'o651;
		14'h2ff: data = 9'o652;
		14'h300: data = 9'o552;
		14'h301: data = 9'o552;
		14'h302: data = 9'o552;
		14'h303: data = 9'o652;
		14'h304: data = 9'o652;
		14'h305: data = 9'o652;
		14'h306: data = 9'o652;
		14'h307: data = 9'o652;
		14'h308: data = 9'o552;
		14'h309: data = 9'o652;
		14'h30a: data = 9'o651;
		14'h30b: data = 9'o651;
		14'h30c: data = 9'o652;
		14'h30d: data = 9'o552;
		14'h30e: data = 9'o551;
		14'h30f: data = 9'o552;
		14'h310: data = 9'o652;
		14'h311: data = 9'o551;
		14'h312: data = 9'o551;
		14'h313: data = 9'o651;
		14'h314: data = 9'o651;
		14'h315: data = 9'o651;
		14'h316: data = 9'o0;
		14'h317: data = 9'o0;
		14'h318: data = 9'o0;
		14'h319: data = 9'o0;
		14'h31a: data = 9'o0;
		14'h31b: data = 9'o0;
		14'h31c: data = 9'o0;
		14'h31d: data = 9'o0;
		14'h31e: data = 9'o0;
		14'h31f: data = 9'o0;
		14'h320: data = 9'o0;
		14'h321: data = 9'o0;
		14'h322: data = 9'o0;
		14'h323: data = 9'o0;
		14'h324: data = 9'o0;
		14'h325: data = 9'o0;
		14'h326: data = 9'o0;
		14'h327: data = 9'o652;
		14'h328: data = 9'o662;
		14'h329: data = 9'o773;
		14'h32a: data = 9'o773;
		14'h32b: data = 9'o773;
		14'h32c: data = 9'o773;
		14'h32d: data = 9'o773;
		14'h32e: data = 9'o773;
		14'h32f: data = 9'o773;
		14'h330: data = 9'o773;
		14'h331: data = 9'o773;
		14'h332: data = 9'o773;
		14'h333: data = 9'o773;
		14'h334: data = 9'o773;
		14'h335: data = 9'o773;
		14'h336: data = 9'o773;
		14'h337: data = 9'o773;
		14'h338: data = 9'o773;
		14'h339: data = 9'o773;
		14'h33a: data = 9'o773;
		14'h33b: data = 9'o773;
		14'h33c: data = 9'o773;
		14'h33d: data = 9'o773;
		14'h33e: data = 9'o773;
		14'h33f: data = 9'o773;
		14'h340: data = 9'o773;
		14'h341: data = 9'o773;
		14'h342: data = 9'o773;
		14'h343: data = 9'o773;
		14'h344: data = 9'o773;
		14'h345: data = 9'o773;
		14'h346: data = 9'o773;
		14'h347: data = 9'o773;
		14'h348: data = 9'o773;
		14'h349: data = 9'o773;
		14'h34a: data = 9'o773;
		14'h34b: data = 9'o773;
		14'h34c: data = 9'o773;
		14'h34d: data = 9'o773;
		14'h34e: data = 9'o773;
		14'h34f: data = 9'o773;
		14'h350: data = 9'o773;
		14'h351: data = 9'o773;
		14'h352: data = 9'o773;
		14'h353: data = 9'o773;
		14'h354: data = 9'o773;
		14'h355: data = 9'o773;
		14'h356: data = 9'o773;
		14'h357: data = 9'o773;
		14'h358: data = 9'o773;
		14'h359: data = 9'o773;
		14'h35a: data = 9'o773;
		14'h35b: data = 9'o773;
		14'h35c: data = 9'o773;
		14'h35d: data = 9'o773;
		14'h35e: data = 9'o773;
		14'h35f: data = 9'o773;
		14'h360: data = 9'o773;
		14'h361: data = 9'o773;
		14'h362: data = 9'o773;
		14'h363: data = 9'o773;
		14'h364: data = 9'o773;
		14'h365: data = 9'o773;
		14'h366: data = 9'o773;
		14'h367: data = 9'o773;
		14'h368: data = 9'o773;
		14'h369: data = 9'o773;
		14'h36a: data = 9'o773;
		14'h36b: data = 9'o773;
		14'h36c: data = 9'o773;
		14'h36d: data = 9'o773;
		14'h36e: data = 9'o773;
		14'h36f: data = 9'o773;
		14'h370: data = 9'o773;
		14'h371: data = 9'o773;
		14'h372: data = 9'o773;
		14'h373: data = 9'o773;
		14'h374: data = 9'o773;
		14'h375: data = 9'o773;
		14'h376: data = 9'o773;
		14'h377: data = 9'o773;
		14'h378: data = 9'o773;
		14'h379: data = 9'o762;
		14'h37a: data = 9'o0;
		14'h37b: data = 9'o0;
		14'h37c: data = 9'o0;
		14'h37d: data = 9'o0;
		14'h37e: data = 9'o0;
		14'h37f: data = 9'o0;
		14'h380: data = 9'o0;
		14'h381: data = 9'o0;
		14'h382: data = 9'o0;
		14'h383: data = 9'o0;
		14'h384: data = 9'o0;
		14'h385: data = 9'o0;
		14'h386: data = 9'o0;
		14'h387: data = 9'o0;
		14'h388: data = 9'o0;
		14'h389: data = 9'o0;
		14'h38a: data = 9'o0;
		14'h38b: data = 9'o551;
		14'h38c: data = 9'o762;
		14'h38d: data = 9'o773;
		14'h38e: data = 9'o773;
		14'h38f: data = 9'o773;
		14'h390: data = 9'o773;
		14'h391: data = 9'o773;
		14'h392: data = 9'o773;
		14'h393: data = 9'o773;
		14'h394: data = 9'o773;
		14'h395: data = 9'o773;
		14'h396: data = 9'o773;
		14'h397: data = 9'o773;
		14'h398: data = 9'o773;
		14'h399: data = 9'o773;
		14'h39a: data = 9'o773;
		14'h39b: data = 9'o773;
		14'h39c: data = 9'o773;
		14'h39d: data = 9'o773;
		14'h39e: data = 9'o773;
		14'h39f: data = 9'o773;
		14'h3a0: data = 9'o773;
		14'h3a1: data = 9'o773;
		14'h3a2: data = 9'o773;
		14'h3a3: data = 9'o773;
		14'h3a4: data = 9'o773;
		14'h3a5: data = 9'o773;
		14'h3a6: data = 9'o773;
		14'h3a7: data = 9'o773;
		14'h3a8: data = 9'o773;
		14'h3a9: data = 9'o773;
		14'h3aa: data = 9'o773;
		14'h3ab: data = 9'o773;
		14'h3ac: data = 9'o773;
		14'h3ad: data = 9'o773;
		14'h3ae: data = 9'o773;
		14'h3af: data = 9'o773;
		14'h3b0: data = 9'o773;
		14'h3b1: data = 9'o773;
		14'h3b2: data = 9'o773;
		14'h3b3: data = 9'o773;
		14'h3b4: data = 9'o773;
		14'h3b5: data = 9'o773;
		14'h3b6: data = 9'o773;
		14'h3b7: data = 9'o773;
		14'h3b8: data = 9'o773;
		14'h3b9: data = 9'o773;
		14'h3ba: data = 9'o773;
		14'h3bb: data = 9'o773;
		14'h3bc: data = 9'o773;
		14'h3bd: data = 9'o773;
		14'h3be: data = 9'o773;
		14'h3bf: data = 9'o773;
		14'h3c0: data = 9'o773;
		14'h3c1: data = 9'o773;
		14'h3c2: data = 9'o773;
		14'h3c3: data = 9'o773;
		14'h3c4: data = 9'o773;
		14'h3c5: data = 9'o773;
		14'h3c6: data = 9'o773;
		14'h3c7: data = 9'o773;
		14'h3c8: data = 9'o773;
		14'h3c9: data = 9'o773;
		14'h3ca: data = 9'o773;
		14'h3cb: data = 9'o773;
		14'h3cc: data = 9'o773;
		14'h3cd: data = 9'o773;
		14'h3ce: data = 9'o773;
		14'h3cf: data = 9'o773;
		14'h3d0: data = 9'o773;
		14'h3d1: data = 9'o773;
		14'h3d2: data = 9'o773;
		14'h3d3: data = 9'o773;
		14'h3d4: data = 9'o773;
		14'h3d5: data = 9'o773;
		14'h3d6: data = 9'o773;
		14'h3d7: data = 9'o773;
		14'h3d8: data = 9'o773;
		14'h3d9: data = 9'o773;
		14'h3da: data = 9'o773;
		14'h3db: data = 9'o773;
		14'h3dc: data = 9'o773;
		14'h3dd: data = 9'o762;
		14'h3de: data = 9'o0;
		14'h3df: data = 9'o0;
		14'h3e0: data = 9'o0;
		14'h3e1: data = 9'o0;
		14'h3e2: data = 9'o0;
		14'h3e3: data = 9'o0;
		14'h3e4: data = 9'o0;
		14'h3e5: data = 9'o0;
		14'h3e6: data = 9'o0;
		14'h3e7: data = 9'o0;
		14'h3e8: data = 9'o0;
		14'h3e9: data = 9'o0;
		14'h3ea: data = 9'o0;
		14'h3eb: data = 9'o0;
		14'h3ec: data = 9'o0;
		14'h3ed: data = 9'o0;
		14'h3ee: data = 9'o0;
		14'h3ef: data = 9'o651;
		14'h3f0: data = 9'o762;
		14'h3f1: data = 9'o773;
		14'h3f2: data = 9'o773;
		14'h3f3: data = 9'o773;
		14'h3f4: data = 9'o773;
		14'h3f5: data = 9'o773;
		14'h3f6: data = 9'o773;
		14'h3f7: data = 9'o773;
		14'h3f8: data = 9'o773;
		14'h3f9: data = 9'o773;
		14'h3fa: data = 9'o773;
		14'h3fb: data = 9'o773;
		14'h3fc: data = 9'o773;
		14'h3fd: data = 9'o773;
		14'h3fe: data = 9'o773;
		14'h3ff: data = 9'o773;
		14'h400: data = 9'o773;
		14'h401: data = 9'o773;
		14'h402: data = 9'o773;
		14'h403: data = 9'o773;
		14'h404: data = 9'o773;
		14'h405: data = 9'o773;
		14'h406: data = 9'o773;
		14'h407: data = 9'o773;
		14'h408: data = 9'o773;
		14'h409: data = 9'o773;
		14'h40a: data = 9'o773;
		14'h40b: data = 9'o773;
		14'h40c: data = 9'o773;
		14'h40d: data = 9'o773;
		14'h40e: data = 9'o773;
		14'h40f: data = 9'o773;
		14'h410: data = 9'o773;
		14'h411: data = 9'o773;
		14'h412: data = 9'o773;
		14'h413: data = 9'o773;
		14'h414: data = 9'o773;
		14'h415: data = 9'o773;
		14'h416: data = 9'o773;
		14'h417: data = 9'o773;
		14'h418: data = 9'o773;
		14'h419: data = 9'o773;
		14'h41a: data = 9'o773;
		14'h41b: data = 9'o773;
		14'h41c: data = 9'o773;
		14'h41d: data = 9'o773;
		14'h41e: data = 9'o773;
		14'h41f: data = 9'o773;
		14'h420: data = 9'o773;
		14'h421: data = 9'o773;
		14'h422: data = 9'o773;
		14'h423: data = 9'o773;
		14'h424: data = 9'o773;
		14'h425: data = 9'o773;
		14'h426: data = 9'o773;
		14'h427: data = 9'o773;
		14'h428: data = 9'o773;
		14'h429: data = 9'o773;
		14'h42a: data = 9'o773;
		14'h42b: data = 9'o773;
		14'h42c: data = 9'o773;
		14'h42d: data = 9'o773;
		14'h42e: data = 9'o773;
		14'h42f: data = 9'o773;
		14'h430: data = 9'o773;
		14'h431: data = 9'o773;
		14'h432: data = 9'o773;
		14'h433: data = 9'o773;
		14'h434: data = 9'o773;
		14'h435: data = 9'o773;
		14'h436: data = 9'o773;
		14'h437: data = 9'o773;
		14'h438: data = 9'o773;
		14'h439: data = 9'o773;
		14'h43a: data = 9'o773;
		14'h43b: data = 9'o773;
		14'h43c: data = 9'o773;
		14'h43d: data = 9'o773;
		14'h43e: data = 9'o773;
		14'h43f: data = 9'o773;
		14'h440: data = 9'o773;
		14'h441: data = 9'o763;
		14'h442: data = 9'o0;
		14'h443: data = 9'o0;
		14'h444: data = 9'o0;
		14'h445: data = 9'o0;
		14'h446: data = 9'o0;
		14'h447: data = 9'o0;
		14'h448: data = 9'o0;
		14'h449: data = 9'o0;
		14'h44a: data = 9'o0;
		14'h44b: data = 9'o0;
		14'h44c: data = 9'o0;
		14'h44d: data = 9'o0;
		14'h44e: data = 9'o0;
		14'h44f: data = 9'o0;
		14'h450: data = 9'o0;
		14'h451: data = 9'o0;
		14'h452: data = 9'o0;
		14'h453: data = 9'o651;
		14'h454: data = 9'o762;
		14'h455: data = 9'o773;
		14'h456: data = 9'o773;
		14'h457: data = 9'o773;
		14'h458: data = 9'o773;
		14'h459: data = 9'o773;
		14'h45a: data = 9'o773;
		14'h45b: data = 9'o773;
		14'h45c: data = 9'o773;
		14'h45d: data = 9'o773;
		14'h45e: data = 9'o773;
		14'h45f: data = 9'o773;
		14'h460: data = 9'o773;
		14'h461: data = 9'o773;
		14'h462: data = 9'o773;
		14'h463: data = 9'o773;
		14'h464: data = 9'o773;
		14'h465: data = 9'o773;
		14'h466: data = 9'o773;
		14'h467: data = 9'o773;
		14'h468: data = 9'o773;
		14'h469: data = 9'o773;
		14'h46a: data = 9'o773;
		14'h46b: data = 9'o773;
		14'h46c: data = 9'o773;
		14'h46d: data = 9'o773;
		14'h46e: data = 9'o773;
		14'h46f: data = 9'o773;
		14'h470: data = 9'o773;
		14'h471: data = 9'o773;
		14'h472: data = 9'o773;
		14'h473: data = 9'o773;
		14'h474: data = 9'o773;
		14'h475: data = 9'o773;
		14'h476: data = 9'o773;
		14'h477: data = 9'o773;
		14'h478: data = 9'o773;
		14'h479: data = 9'o773;
		14'h47a: data = 9'o773;
		14'h47b: data = 9'o773;
		14'h47c: data = 9'o773;
		14'h47d: data = 9'o773;
		14'h47e: data = 9'o773;
		14'h47f: data = 9'o773;
		14'h480: data = 9'o773;
		14'h481: data = 9'o773;
		14'h482: data = 9'o773;
		14'h483: data = 9'o773;
		14'h484: data = 9'o773;
		14'h485: data = 9'o773;
		14'h486: data = 9'o773;
		14'h487: data = 9'o773;
		14'h488: data = 9'o773;
		14'h489: data = 9'o773;
		14'h48a: data = 9'o773;
		14'h48b: data = 9'o773;
		14'h48c: data = 9'o773;
		14'h48d: data = 9'o773;
		14'h48e: data = 9'o773;
		14'h48f: data = 9'o773;
		14'h490: data = 9'o773;
		14'h491: data = 9'o773;
		14'h492: data = 9'o773;
		14'h493: data = 9'o773;
		14'h494: data = 9'o773;
		14'h495: data = 9'o773;
		14'h496: data = 9'o773;
		14'h497: data = 9'o773;
		14'h498: data = 9'o773;
		14'h499: data = 9'o773;
		14'h49a: data = 9'o773;
		14'h49b: data = 9'o773;
		14'h49c: data = 9'o773;
		14'h49d: data = 9'o773;
		14'h49e: data = 9'o773;
		14'h49f: data = 9'o773;
		14'h4a0: data = 9'o773;
		14'h4a1: data = 9'o773;
		14'h4a2: data = 9'o773;
		14'h4a3: data = 9'o773;
		14'h4a4: data = 9'o773;
		14'h4a5: data = 9'o763;
		14'h4a6: data = 9'o0;
		14'h4a7: data = 9'o0;
		14'h4a8: data = 9'o0;
		14'h4a9: data = 9'o0;
		14'h4aa: data = 9'o0;
		14'h4ab: data = 9'o0;
		14'h4ac: data = 9'o0;
		14'h4ad: data = 9'o0;
		14'h4ae: data = 9'o0;
		14'h4af: data = 9'o0;
		14'h4b0: data = 9'o0;
		14'h4b1: data = 9'o0;
		14'h4b2: data = 9'o0;
		14'h4b3: data = 9'o0;
		14'h4b4: data = 9'o0;
		14'h4b5: data = 9'o0;
		14'h4b6: data = 9'o0;
		14'h4b7: data = 9'o651;
		14'h4b8: data = 9'o762;
		14'h4b9: data = 9'o773;
		14'h4ba: data = 9'o773;
		14'h4bb: data = 9'o773;
		14'h4bc: data = 9'o773;
		14'h4bd: data = 9'o773;
		14'h4be: data = 9'o773;
		14'h4bf: data = 9'o773;
		14'h4c0: data = 9'o773;
		14'h4c1: data = 9'o773;
		14'h4c2: data = 9'o773;
		14'h4c3: data = 9'o773;
		14'h4c4: data = 9'o773;
		14'h4c5: data = 9'o773;
		14'h4c6: data = 9'o773;
		14'h4c7: data = 9'o773;
		14'h4c8: data = 9'o773;
		14'h4c9: data = 9'o773;
		14'h4ca: data = 9'o773;
		14'h4cb: data = 9'o773;
		14'h4cc: data = 9'o773;
		14'h4cd: data = 9'o773;
		14'h4ce: data = 9'o773;
		14'h4cf: data = 9'o773;
		14'h4d0: data = 9'o773;
		14'h4d1: data = 9'o773;
		14'h4d2: data = 9'o773;
		14'h4d3: data = 9'o773;
		14'h4d4: data = 9'o773;
		14'h4d5: data = 9'o773;
		14'h4d6: data = 9'o773;
		14'h4d7: data = 9'o773;
		14'h4d8: data = 9'o773;
		14'h4d9: data = 9'o773;
		14'h4da: data = 9'o773;
		14'h4db: data = 9'o773;
		14'h4dc: data = 9'o773;
		14'h4dd: data = 9'o773;
		14'h4de: data = 9'o773;
		14'h4df: data = 9'o773;
		14'h4e0: data = 9'o773;
		14'h4e1: data = 9'o773;
		14'h4e2: data = 9'o773;
		14'h4e3: data = 9'o773;
		14'h4e4: data = 9'o773;
		14'h4e5: data = 9'o773;
		14'h4e6: data = 9'o773;
		14'h4e7: data = 9'o773;
		14'h4e8: data = 9'o773;
		14'h4e9: data = 9'o773;
		14'h4ea: data = 9'o773;
		14'h4eb: data = 9'o773;
		14'h4ec: data = 9'o773;
		14'h4ed: data = 9'o773;
		14'h4ee: data = 9'o773;
		14'h4ef: data = 9'o773;
		14'h4f0: data = 9'o773;
		14'h4f1: data = 9'o773;
		14'h4f2: data = 9'o773;
		14'h4f3: data = 9'o773;
		14'h4f4: data = 9'o773;
		14'h4f5: data = 9'o773;
		14'h4f6: data = 9'o773;
		14'h4f7: data = 9'o773;
		14'h4f8: data = 9'o773;
		14'h4f9: data = 9'o773;
		14'h4fa: data = 9'o773;
		14'h4fb: data = 9'o773;
		14'h4fc: data = 9'o773;
		14'h4fd: data = 9'o773;
		14'h4fe: data = 9'o773;
		14'h4ff: data = 9'o773;
		14'h500: data = 9'o773;
		14'h501: data = 9'o773;
		14'h502: data = 9'o773;
		14'h503: data = 9'o773;
		14'h504: data = 9'o773;
		14'h505: data = 9'o773;
		14'h506: data = 9'o773;
		14'h507: data = 9'o773;
		14'h508: data = 9'o773;
		14'h509: data = 9'o762;
		14'h50a: data = 9'o0;
		14'h50b: data = 9'o0;
		14'h50c: data = 9'o0;
		14'h50d: data = 9'o0;
		14'h50e: data = 9'o0;
		14'h50f: data = 9'o0;
		14'h510: data = 9'o0;
		14'h511: data = 9'o0;
		14'h512: data = 9'o0;
		14'h513: data = 9'o0;
		14'h514: data = 9'o0;
		14'h515: data = 9'o0;
		14'h516: data = 9'o0;
		14'h517: data = 9'o0;
		14'h518: data = 9'o0;
		14'h519: data = 9'o0;
		14'h51a: data = 9'o0;
		14'h51b: data = 9'o651;
		14'h51c: data = 9'o762;
		14'h51d: data = 9'o773;
		14'h51e: data = 9'o773;
		14'h51f: data = 9'o773;
		14'h520: data = 9'o773;
		14'h521: data = 9'o773;
		14'h522: data = 9'o773;
		14'h523: data = 9'o773;
		14'h524: data = 9'o773;
		14'h525: data = 9'o773;
		14'h526: data = 9'o773;
		14'h527: data = 9'o773;
		14'h528: data = 9'o773;
		14'h529: data = 9'o773;
		14'h52a: data = 9'o773;
		14'h52b: data = 9'o773;
		14'h52c: data = 9'o773;
		14'h52d: data = 9'o773;
		14'h52e: data = 9'o773;
		14'h52f: data = 9'o773;
		14'h530: data = 9'o773;
		14'h531: data = 9'o773;
		14'h532: data = 9'o773;
		14'h533: data = 9'o773;
		14'h534: data = 9'o773;
		14'h535: data = 9'o773;
		14'h536: data = 9'o773;
		14'h537: data = 9'o773;
		14'h538: data = 9'o773;
		14'h539: data = 9'o773;
		14'h53a: data = 9'o773;
		14'h53b: data = 9'o773;
		14'h53c: data = 9'o773;
		14'h53d: data = 9'o773;
		14'h53e: data = 9'o773;
		14'h53f: data = 9'o773;
		14'h540: data = 9'o773;
		14'h541: data = 9'o773;
		14'h542: data = 9'o773;
		14'h543: data = 9'o773;
		14'h544: data = 9'o773;
		14'h545: data = 9'o773;
		14'h546: data = 9'o773;
		14'h547: data = 9'o773;
		14'h548: data = 9'o773;
		14'h549: data = 9'o773;
		14'h54a: data = 9'o773;
		14'h54b: data = 9'o773;
		14'h54c: data = 9'o773;
		14'h54d: data = 9'o773;
		14'h54e: data = 9'o773;
		14'h54f: data = 9'o773;
		14'h550: data = 9'o773;
		14'h551: data = 9'o773;
		14'h552: data = 9'o773;
		14'h553: data = 9'o773;
		14'h554: data = 9'o773;
		14'h555: data = 9'o773;
		14'h556: data = 9'o773;
		14'h557: data = 9'o773;
		14'h558: data = 9'o773;
		14'h559: data = 9'o773;
		14'h55a: data = 9'o773;
		14'h55b: data = 9'o773;
		14'h55c: data = 9'o773;
		14'h55d: data = 9'o773;
		14'h55e: data = 9'o773;
		14'h55f: data = 9'o773;
		14'h560: data = 9'o773;
		14'h561: data = 9'o773;
		14'h562: data = 9'o773;
		14'h563: data = 9'o773;
		14'h564: data = 9'o773;
		14'h565: data = 9'o773;
		14'h566: data = 9'o773;
		14'h567: data = 9'o773;
		14'h568: data = 9'o773;
		14'h569: data = 9'o773;
		14'h56a: data = 9'o773;
		14'h56b: data = 9'o773;
		14'h56c: data = 9'o773;
		14'h56d: data = 9'o762;
		14'h56e: data = 9'o0;
		14'h56f: data = 9'o0;
		14'h570: data = 9'o0;
		14'h571: data = 9'o0;
		14'h572: data = 9'o0;
		14'h573: data = 9'o0;
		14'h574: data = 9'o0;
		14'h575: data = 9'o0;
		14'h576: data = 9'o0;
		14'h577: data = 9'o0;
		14'h578: data = 9'o0;
		14'h579: data = 9'o0;
		14'h57a: data = 9'o0;
		14'h57b: data = 9'o0;
		14'h57c: data = 9'o0;
		14'h57d: data = 9'o0;
		14'h57e: data = 9'o0;
		14'h57f: data = 9'o651;
		14'h580: data = 9'o762;
		14'h581: data = 9'o773;
		14'h582: data = 9'o773;
		14'h583: data = 9'o773;
		14'h584: data = 9'o773;
		14'h585: data = 9'o773;
		14'h586: data = 9'o773;
		14'h587: data = 9'o773;
		14'h588: data = 9'o773;
		14'h589: data = 9'o773;
		14'h58a: data = 9'o773;
		14'h58b: data = 9'o773;
		14'h58c: data = 9'o773;
		14'h58d: data = 9'o773;
		14'h58e: data = 9'o773;
		14'h58f: data = 9'o773;
		14'h590: data = 9'o773;
		14'h591: data = 9'o773;
		14'h592: data = 9'o773;
		14'h593: data = 9'o773;
		14'h594: data = 9'o773;
		14'h595: data = 9'o773;
		14'h596: data = 9'o773;
		14'h597: data = 9'o773;
		14'h598: data = 9'o773;
		14'h599: data = 9'o773;
		14'h59a: data = 9'o773;
		14'h59b: data = 9'o773;
		14'h59c: data = 9'o773;
		14'h59d: data = 9'o773;
		14'h59e: data = 9'o773;
		14'h59f: data = 9'o773;
		14'h5a0: data = 9'o773;
		14'h5a1: data = 9'o773;
		14'h5a2: data = 9'o773;
		14'h5a3: data = 9'o773;
		14'h5a4: data = 9'o773;
		14'h5a5: data = 9'o773;
		14'h5a6: data = 9'o773;
		14'h5a7: data = 9'o773;
		14'h5a8: data = 9'o773;
		14'h5a9: data = 9'o773;
		14'h5aa: data = 9'o773;
		14'h5ab: data = 9'o773;
		14'h5ac: data = 9'o773;
		14'h5ad: data = 9'o773;
		14'h5ae: data = 9'o773;
		14'h5af: data = 9'o773;
		14'h5b0: data = 9'o773;
		14'h5b1: data = 9'o773;
		14'h5b2: data = 9'o773;
		14'h5b3: data = 9'o773;
		14'h5b4: data = 9'o773;
		14'h5b5: data = 9'o773;
		14'h5b6: data = 9'o773;
		14'h5b7: data = 9'o773;
		14'h5b8: data = 9'o773;
		14'h5b9: data = 9'o773;
		14'h5ba: data = 9'o773;
		14'h5bb: data = 9'o773;
		14'h5bc: data = 9'o773;
		14'h5bd: data = 9'o773;
		14'h5be: data = 9'o773;
		14'h5bf: data = 9'o773;
		14'h5c0: data = 9'o773;
		14'h5c1: data = 9'o773;
		14'h5c2: data = 9'o773;
		14'h5c3: data = 9'o773;
		14'h5c4: data = 9'o773;
		14'h5c5: data = 9'o773;
		14'h5c6: data = 9'o773;
		14'h5c7: data = 9'o773;
		14'h5c8: data = 9'o773;
		14'h5c9: data = 9'o773;
		14'h5ca: data = 9'o773;
		14'h5cb: data = 9'o773;
		14'h5cc: data = 9'o773;
		14'h5cd: data = 9'o773;
		14'h5ce: data = 9'o773;
		14'h5cf: data = 9'o773;
		14'h5d0: data = 9'o773;
		14'h5d1: data = 9'o763;
		14'h5d2: data = 9'o0;
		14'h5d3: data = 9'o0;
		14'h5d4: data = 9'o0;
		14'h5d5: data = 9'o0;
		14'h5d6: data = 9'o0;
		14'h5d7: data = 9'o0;
		14'h5d8: data = 9'o0;
		14'h5d9: data = 9'o0;
		14'h5da: data = 9'o0;
		14'h5db: data = 9'o0;
		14'h5dc: data = 9'o0;
		14'h5dd: data = 9'o0;
		14'h5de: data = 9'o0;
		14'h5df: data = 9'o0;
		14'h5e0: data = 9'o0;
		14'h5e1: data = 9'o0;
		14'h5e2: data = 9'o0;
		14'h5e3: data = 9'o651;
		14'h5e4: data = 9'o762;
		14'h5e5: data = 9'o773;
		14'h5e6: data = 9'o773;
		14'h5e7: data = 9'o773;
		14'h5e8: data = 9'o773;
		14'h5e9: data = 9'o773;
		14'h5ea: data = 9'o773;
		14'h5eb: data = 9'o773;
		14'h5ec: data = 9'o773;
		14'h5ed: data = 9'o773;
		14'h5ee: data = 9'o773;
		14'h5ef: data = 9'o773;
		14'h5f0: data = 9'o773;
		14'h5f1: data = 9'o773;
		14'h5f2: data = 9'o773;
		14'h5f3: data = 9'o773;
		14'h5f4: data = 9'o773;
		14'h5f5: data = 9'o773;
		14'h5f6: data = 9'o773;
		14'h5f7: data = 9'o773;
		14'h5f8: data = 9'o773;
		14'h5f9: data = 9'o773;
		14'h5fa: data = 9'o773;
		14'h5fb: data = 9'o773;
		14'h5fc: data = 9'o773;
		14'h5fd: data = 9'o773;
		14'h5fe: data = 9'o773;
		14'h5ff: data = 9'o773;
		14'h600: data = 9'o773;
		14'h601: data = 9'o773;
		14'h602: data = 9'o773;
		14'h603: data = 9'o773;
		14'h604: data = 9'o773;
		14'h605: data = 9'o773;
		14'h606: data = 9'o773;
		14'h607: data = 9'o773;
		14'h608: data = 9'o773;
		14'h609: data = 9'o773;
		14'h60a: data = 9'o773;
		14'h60b: data = 9'o773;
		14'h60c: data = 9'o773;
		14'h60d: data = 9'o773;
		14'h60e: data = 9'o773;
		14'h60f: data = 9'o773;
		14'h610: data = 9'o773;
		14'h611: data = 9'o773;
		14'h612: data = 9'o773;
		14'h613: data = 9'o773;
		14'h614: data = 9'o773;
		14'h615: data = 9'o773;
		14'h616: data = 9'o773;
		14'h617: data = 9'o773;
		14'h618: data = 9'o773;
		14'h619: data = 9'o773;
		14'h61a: data = 9'o773;
		14'h61b: data = 9'o773;
		14'h61c: data = 9'o773;
		14'h61d: data = 9'o773;
		14'h61e: data = 9'o773;
		14'h61f: data = 9'o773;
		14'h620: data = 9'o773;
		14'h621: data = 9'o773;
		14'h622: data = 9'o773;
		14'h623: data = 9'o773;
		14'h624: data = 9'o773;
		14'h625: data = 9'o773;
		14'h626: data = 9'o773;
		14'h627: data = 9'o773;
		14'h628: data = 9'o773;
		14'h629: data = 9'o773;
		14'h62a: data = 9'o773;
		14'h62b: data = 9'o773;
		14'h62c: data = 9'o773;
		14'h62d: data = 9'o773;
		14'h62e: data = 9'o773;
		14'h62f: data = 9'o773;
		14'h630: data = 9'o773;
		14'h631: data = 9'o773;
		14'h632: data = 9'o773;
		14'h633: data = 9'o773;
		14'h634: data = 9'o773;
		14'h635: data = 9'o763;
		14'h636: data = 9'o0;
		14'h637: data = 9'o0;
		14'h638: data = 9'o0;
		14'h639: data = 9'o0;
		14'h63a: data = 9'o0;
		14'h63b: data = 9'o0;
		14'h63c: data = 9'o0;
		14'h63d: data = 9'o0;
		14'h63e: data = 9'o0;
		14'h63f: data = 9'o0;
		14'h640: data = 9'o0;
		14'h641: data = 9'o0;
		14'h642: data = 9'o0;
		14'h643: data = 9'o0;
		14'h644: data = 9'o0;
		14'h645: data = 9'o0;
		14'h646: data = 9'o0;
		14'h647: data = 9'o651;
		14'h648: data = 9'o762;
		14'h649: data = 9'o773;
		14'h64a: data = 9'o773;
		14'h64b: data = 9'o773;
		14'h64c: data = 9'o773;
		14'h64d: data = 9'o773;
		14'h64e: data = 9'o773;
		14'h64f: data = 9'o773;
		14'h650: data = 9'o773;
		14'h651: data = 9'o773;
		14'h652: data = 9'o773;
		14'h653: data = 9'o773;
		14'h654: data = 9'o773;
		14'h655: data = 9'o773;
		14'h656: data = 9'o773;
		14'h657: data = 9'o773;
		14'h658: data = 9'o773;
		14'h659: data = 9'o773;
		14'h65a: data = 9'o773;
		14'h65b: data = 9'o773;
		14'h65c: data = 9'o773;
		14'h65d: data = 9'o773;
		14'h65e: data = 9'o773;
		14'h65f: data = 9'o773;
		14'h660: data = 9'o773;
		14'h661: data = 9'o773;
		14'h662: data = 9'o773;
		14'h663: data = 9'o773;
		14'h664: data = 9'o773;
		14'h665: data = 9'o773;
		14'h666: data = 9'o773;
		14'h667: data = 9'o773;
		14'h668: data = 9'o773;
		14'h669: data = 9'o773;
		14'h66a: data = 9'o773;
		14'h66b: data = 9'o773;
		14'h66c: data = 9'o773;
		14'h66d: data = 9'o773;
		14'h66e: data = 9'o773;
		14'h66f: data = 9'o773;
		14'h670: data = 9'o773;
		14'h671: data = 9'o773;
		14'h672: data = 9'o773;
		14'h673: data = 9'o773;
		14'h674: data = 9'o773;
		14'h675: data = 9'o773;
		14'h676: data = 9'o773;
		14'h677: data = 9'o773;
		14'h678: data = 9'o773;
		14'h679: data = 9'o773;
		14'h67a: data = 9'o773;
		14'h67b: data = 9'o773;
		14'h67c: data = 9'o773;
		14'h67d: data = 9'o773;
		14'h67e: data = 9'o773;
		14'h67f: data = 9'o773;
		14'h680: data = 9'o773;
		14'h681: data = 9'o773;
		14'h682: data = 9'o773;
		14'h683: data = 9'o773;
		14'h684: data = 9'o773;
		14'h685: data = 9'o773;
		14'h686: data = 9'o773;
		14'h687: data = 9'o773;
		14'h688: data = 9'o773;
		14'h689: data = 9'o773;
		14'h68a: data = 9'o773;
		14'h68b: data = 9'o773;
		14'h68c: data = 9'o773;
		14'h68d: data = 9'o773;
		14'h68e: data = 9'o773;
		14'h68f: data = 9'o773;
		14'h690: data = 9'o773;
		14'h691: data = 9'o773;
		14'h692: data = 9'o773;
		14'h693: data = 9'o773;
		14'h694: data = 9'o773;
		14'h695: data = 9'o773;
		14'h696: data = 9'o773;
		14'h697: data = 9'o773;
		14'h698: data = 9'o773;
		14'h699: data = 9'o762;
		14'h69a: data = 9'o0;
		14'h69b: data = 9'o0;
		14'h69c: data = 9'o0;
		14'h69d: data = 9'o0;
		14'h69e: data = 9'o0;
		14'h69f: data = 9'o0;
		14'h6a0: data = 9'o0;
		14'h6a1: data = 9'o0;
		14'h6a2: data = 9'o0;
		14'h6a3: data = 9'o0;
		14'h6a4: data = 9'o0;
		14'h6a5: data = 9'o0;
		14'h6a6: data = 9'o0;
		14'h6a7: data = 9'o0;
		14'h6a8: data = 9'o0;
		14'h6a9: data = 9'o0;
		14'h6aa: data = 9'o0;
		14'h6ab: data = 9'o651;
		14'h6ac: data = 9'o762;
		14'h6ad: data = 9'o773;
		14'h6ae: data = 9'o773;
		14'h6af: data = 9'o773;
		14'h6b0: data = 9'o773;
		14'h6b1: data = 9'o773;
		14'h6b2: data = 9'o773;
		14'h6b3: data = 9'o773;
		14'h6b4: data = 9'o773;
		14'h6b5: data = 9'o773;
		14'h6b6: data = 9'o773;
		14'h6b7: data = 9'o773;
		14'h6b8: data = 9'o773;
		14'h6b9: data = 9'o773;
		14'h6ba: data = 9'o773;
		14'h6bb: data = 9'o773;
		14'h6bc: data = 9'o773;
		14'h6bd: data = 9'o773;
		14'h6be: data = 9'o773;
		14'h6bf: data = 9'o773;
		14'h6c0: data = 9'o773;
		14'h6c1: data = 9'o773;
		14'h6c2: data = 9'o773;
		14'h6c3: data = 9'o773;
		14'h6c4: data = 9'o773;
		14'h6c5: data = 9'o773;
		14'h6c6: data = 9'o773;
		14'h6c7: data = 9'o773;
		14'h6c8: data = 9'o773;
		14'h6c9: data = 9'o773;
		14'h6ca: data = 9'o773;
		14'h6cb: data = 9'o773;
		14'h6cc: data = 9'o773;
		14'h6cd: data = 9'o773;
		14'h6ce: data = 9'o773;
		14'h6cf: data = 9'o773;
		14'h6d0: data = 9'o773;
		14'h6d1: data = 9'o773;
		14'h6d2: data = 9'o773;
		14'h6d3: data = 9'o773;
		14'h6d4: data = 9'o773;
		14'h6d5: data = 9'o773;
		14'h6d6: data = 9'o773;
		14'h6d7: data = 9'o773;
		14'h6d8: data = 9'o773;
		14'h6d9: data = 9'o773;
		14'h6da: data = 9'o773;
		14'h6db: data = 9'o773;
		14'h6dc: data = 9'o773;
		14'h6dd: data = 9'o773;
		14'h6de: data = 9'o773;
		14'h6df: data = 9'o773;
		14'h6e0: data = 9'o773;
		14'h6e1: data = 9'o773;
		14'h6e2: data = 9'o773;
		14'h6e3: data = 9'o773;
		14'h6e4: data = 9'o773;
		14'h6e5: data = 9'o773;
		14'h6e6: data = 9'o773;
		14'h6e7: data = 9'o773;
		14'h6e8: data = 9'o773;
		14'h6e9: data = 9'o773;
		14'h6ea: data = 9'o773;
		14'h6eb: data = 9'o773;
		14'h6ec: data = 9'o773;
		14'h6ed: data = 9'o773;
		14'h6ee: data = 9'o773;
		14'h6ef: data = 9'o773;
		14'h6f0: data = 9'o773;
		14'h6f1: data = 9'o773;
		14'h6f2: data = 9'o773;
		14'h6f3: data = 9'o773;
		14'h6f4: data = 9'o773;
		14'h6f5: data = 9'o773;
		14'h6f6: data = 9'o773;
		14'h6f7: data = 9'o773;
		14'h6f8: data = 9'o773;
		14'h6f9: data = 9'o773;
		14'h6fa: data = 9'o773;
		14'h6fb: data = 9'o773;
		14'h6fc: data = 9'o773;
		14'h6fd: data = 9'o662;
		14'h6fe: data = 9'o0;
		14'h6ff: data = 9'o0;
		14'h700: data = 9'o0;
		14'h701: data = 9'o0;
		14'h702: data = 9'o0;
		14'h703: data = 9'o0;
		14'h704: data = 9'o0;
		14'h705: data = 9'o0;
		14'h706: data = 9'o0;
		14'h707: data = 9'o0;
		14'h708: data = 9'o0;
		14'h709: data = 9'o0;
		14'h70a: data = 9'o0;
		14'h70b: data = 9'o0;
		14'h70c: data = 9'o0;
		14'h70d: data = 9'o0;
		14'h70e: data = 9'o0;
		14'h70f: data = 9'o651;
		14'h710: data = 9'o762;
		14'h711: data = 9'o773;
		14'h712: data = 9'o773;
		14'h713: data = 9'o773;
		14'h714: data = 9'o773;
		14'h715: data = 9'o773;
		14'h716: data = 9'o773;
		14'h717: data = 9'o773;
		14'h718: data = 9'o773;
		14'h719: data = 9'o773;
		14'h71a: data = 9'o773;
		14'h71b: data = 9'o773;
		14'h71c: data = 9'o773;
		14'h71d: data = 9'o773;
		14'h71e: data = 9'o773;
		14'h71f: data = 9'o773;
		14'h720: data = 9'o773;
		14'h721: data = 9'o773;
		14'h722: data = 9'o773;
		14'h723: data = 9'o773;
		14'h724: data = 9'o773;
		14'h725: data = 9'o773;
		14'h726: data = 9'o773;
		14'h727: data = 9'o773;
		14'h728: data = 9'o773;
		14'h729: data = 9'o773;
		14'h72a: data = 9'o773;
		14'h72b: data = 9'o773;
		14'h72c: data = 9'o773;
		14'h72d: data = 9'o773;
		14'h72e: data = 9'o773;
		14'h72f: data = 9'o773;
		14'h730: data = 9'o773;
		14'h731: data = 9'o773;
		14'h732: data = 9'o773;
		14'h733: data = 9'o773;
		14'h734: data = 9'o773;
		14'h735: data = 9'o773;
		14'h736: data = 9'o773;
		14'h737: data = 9'o773;
		14'h738: data = 9'o673;
		14'h739: data = 9'o673;
		14'h73a: data = 9'o773;
		14'h73b: data = 9'o773;
		14'h73c: data = 9'o773;
		14'h73d: data = 9'o773;
		14'h73e: data = 9'o773;
		14'h73f: data = 9'o773;
		14'h740: data = 9'o773;
		14'h741: data = 9'o773;
		14'h742: data = 9'o773;
		14'h743: data = 9'o773;
		14'h744: data = 9'o773;
		14'h745: data = 9'o773;
		14'h746: data = 9'o773;
		14'h747: data = 9'o773;
		14'h748: data = 9'o773;
		14'h749: data = 9'o773;
		14'h74a: data = 9'o773;
		14'h74b: data = 9'o773;
		14'h74c: data = 9'o773;
		14'h74d: data = 9'o773;
		14'h74e: data = 9'o773;
		14'h74f: data = 9'o773;
		14'h750: data = 9'o773;
		14'h751: data = 9'o773;
		14'h752: data = 9'o773;
		14'h753: data = 9'o773;
		14'h754: data = 9'o773;
		14'h755: data = 9'o773;
		14'h756: data = 9'o773;
		14'h757: data = 9'o773;
		14'h758: data = 9'o773;
		14'h759: data = 9'o773;
		14'h75a: data = 9'o773;
		14'h75b: data = 9'o773;
		14'h75c: data = 9'o773;
		14'h75d: data = 9'o773;
		14'h75e: data = 9'o773;
		14'h75f: data = 9'o773;
		14'h760: data = 9'o773;
		14'h761: data = 9'o762;
		14'h762: data = 9'o0;
		14'h763: data = 9'o0;
		14'h764: data = 9'o0;
		14'h765: data = 9'o0;
		14'h766: data = 9'o0;
		14'h767: data = 9'o0;
		14'h768: data = 9'o0;
		14'h769: data = 9'o0;
		14'h76a: data = 9'o0;
		14'h76b: data = 9'o0;
		14'h76c: data = 9'o0;
		14'h76d: data = 9'o0;
		14'h76e: data = 9'o0;
		14'h76f: data = 9'o0;
		14'h770: data = 9'o0;
		14'h771: data = 9'o0;
		14'h772: data = 9'o0;
		14'h773: data = 9'o651;
		14'h774: data = 9'o762;
		14'h775: data = 9'o773;
		14'h776: data = 9'o773;
		14'h777: data = 9'o773;
		14'h778: data = 9'o773;
		14'h779: data = 9'o773;
		14'h77a: data = 9'o773;
		14'h77b: data = 9'o773;
		14'h77c: data = 9'o773;
		14'h77d: data = 9'o773;
		14'h77e: data = 9'o773;
		14'h77f: data = 9'o773;
		14'h780: data = 9'o773;
		14'h781: data = 9'o773;
		14'h782: data = 9'o773;
		14'h783: data = 9'o773;
		14'h784: data = 9'o773;
		14'h785: data = 9'o773;
		14'h786: data = 9'o773;
		14'h787: data = 9'o773;
		14'h788: data = 9'o773;
		14'h789: data = 9'o773;
		14'h78a: data = 9'o773;
		14'h78b: data = 9'o773;
		14'h78c: data = 9'o773;
		14'h78d: data = 9'o773;
		14'h78e: data = 9'o773;
		14'h78f: data = 9'o773;
		14'h790: data = 9'o773;
		14'h791: data = 9'o773;
		14'h792: data = 9'o773;
		14'h793: data = 9'o773;
		14'h794: data = 9'o773;
		14'h795: data = 9'o773;
		14'h796: data = 9'o773;
		14'h797: data = 9'o773;
		14'h798: data = 9'o773;
		14'h799: data = 9'o773;
		14'h79a: data = 9'o773;
		14'h79b: data = 9'o773;
		14'h79c: data = 9'o573;
		14'h79d: data = 9'o573;
		14'h79e: data = 9'o773;
		14'h79f: data = 9'o773;
		14'h7a0: data = 9'o773;
		14'h7a1: data = 9'o773;
		14'h7a2: data = 9'o773;
		14'h7a3: data = 9'o773;
		14'h7a4: data = 9'o773;
		14'h7a5: data = 9'o773;
		14'h7a6: data = 9'o773;
		14'h7a7: data = 9'o773;
		14'h7a8: data = 9'o773;
		14'h7a9: data = 9'o773;
		14'h7aa: data = 9'o773;
		14'h7ab: data = 9'o773;
		14'h7ac: data = 9'o773;
		14'h7ad: data = 9'o773;
		14'h7ae: data = 9'o773;
		14'h7af: data = 9'o773;
		14'h7b0: data = 9'o773;
		14'h7b1: data = 9'o773;
		14'h7b2: data = 9'o773;
		14'h7b3: data = 9'o773;
		14'h7b4: data = 9'o773;
		14'h7b5: data = 9'o773;
		14'h7b6: data = 9'o773;
		14'h7b7: data = 9'o773;
		14'h7b8: data = 9'o773;
		14'h7b9: data = 9'o773;
		14'h7ba: data = 9'o773;
		14'h7bb: data = 9'o773;
		14'h7bc: data = 9'o773;
		14'h7bd: data = 9'o773;
		14'h7be: data = 9'o773;
		14'h7bf: data = 9'o773;
		14'h7c0: data = 9'o773;
		14'h7c1: data = 9'o773;
		14'h7c2: data = 9'o773;
		14'h7c3: data = 9'o773;
		14'h7c4: data = 9'o773;
		14'h7c5: data = 9'o763;
		14'h7c6: data = 9'o0;
		14'h7c7: data = 9'o0;
		14'h7c8: data = 9'o0;
		14'h7c9: data = 9'o0;
		14'h7ca: data = 9'o0;
		14'h7cb: data = 9'o0;
		14'h7cc: data = 9'o0;
		14'h7cd: data = 9'o0;
		14'h7ce: data = 9'o0;
		14'h7cf: data = 9'o0;
		14'h7d0: data = 9'o0;
		14'h7d1: data = 9'o0;
		14'h7d2: data = 9'o0;
		14'h7d3: data = 9'o0;
		14'h7d4: data = 9'o0;
		14'h7d5: data = 9'o0;
		14'h7d6: data = 9'o0;
		14'h7d7: data = 9'o651;
		14'h7d8: data = 9'o762;
		14'h7d9: data = 9'o773;
		14'h7da: data = 9'o773;
		14'h7db: data = 9'o773;
		14'h7dc: data = 9'o773;
		14'h7dd: data = 9'o773;
		14'h7de: data = 9'o773;
		14'h7df: data = 9'o773;
		14'h7e0: data = 9'o773;
		14'h7e1: data = 9'o773;
		14'h7e2: data = 9'o773;
		14'h7e3: data = 9'o773;
		14'h7e4: data = 9'o773;
		14'h7e5: data = 9'o773;
		14'h7e6: data = 9'o773;
		14'h7e7: data = 9'o773;
		14'h7e8: data = 9'o773;
		14'h7e9: data = 9'o773;
		14'h7ea: data = 9'o773;
		14'h7eb: data = 9'o773;
		14'h7ec: data = 9'o773;
		14'h7ed: data = 9'o773;
		14'h7ee: data = 9'o773;
		14'h7ef: data = 9'o773;
		14'h7f0: data = 9'o773;
		14'h7f1: data = 9'o773;
		14'h7f2: data = 9'o773;
		14'h7f3: data = 9'o773;
		14'h7f4: data = 9'o773;
		14'h7f5: data = 9'o773;
		14'h7f6: data = 9'o773;
		14'h7f7: data = 9'o773;
		14'h7f8: data = 9'o773;
		14'h7f9: data = 9'o773;
		14'h7fa: data = 9'o773;
		14'h7fb: data = 9'o773;
		14'h7fc: data = 9'o773;
		14'h7fd: data = 9'o773;
		14'h7fe: data = 9'o773;
		14'h7ff: data = 9'o773;
		14'h800: data = 9'o463;
		14'h801: data = 9'o362;
		14'h802: data = 9'o773;
		14'h803: data = 9'o773;
		14'h804: data = 9'o773;
		14'h805: data = 9'o773;
		14'h806: data = 9'o773;
		14'h807: data = 9'o773;
		14'h808: data = 9'o773;
		14'h809: data = 9'o773;
		14'h80a: data = 9'o773;
		14'h80b: data = 9'o773;
		14'h80c: data = 9'o773;
		14'h80d: data = 9'o773;
		14'h80e: data = 9'o773;
		14'h80f: data = 9'o773;
		14'h810: data = 9'o773;
		14'h811: data = 9'o773;
		14'h812: data = 9'o773;
		14'h813: data = 9'o773;
		14'h814: data = 9'o773;
		14'h815: data = 9'o773;
		14'h816: data = 9'o773;
		14'h817: data = 9'o773;
		14'h818: data = 9'o773;
		14'h819: data = 9'o773;
		14'h81a: data = 9'o773;
		14'h81b: data = 9'o773;
		14'h81c: data = 9'o773;
		14'h81d: data = 9'o773;
		14'h81e: data = 9'o773;
		14'h81f: data = 9'o773;
		14'h820: data = 9'o773;
		14'h821: data = 9'o773;
		14'h822: data = 9'o773;
		14'h823: data = 9'o773;
		14'h824: data = 9'o773;
		14'h825: data = 9'o773;
		14'h826: data = 9'o773;
		14'h827: data = 9'o773;
		14'h828: data = 9'o773;
		14'h829: data = 9'o763;
		14'h82a: data = 9'o0;
		14'h82b: data = 9'o0;
		14'h82c: data = 9'o0;
		14'h82d: data = 9'o0;
		14'h82e: data = 9'o0;
		14'h82f: data = 9'o0;
		14'h830: data = 9'o0;
		14'h831: data = 9'o0;
		14'h832: data = 9'o0;
		14'h833: data = 9'o0;
		14'h834: data = 9'o0;
		14'h835: data = 9'o0;
		14'h836: data = 9'o0;
		14'h837: data = 9'o0;
		14'h838: data = 9'o0;
		14'h839: data = 9'o0;
		14'h83a: data = 9'o0;
		14'h83b: data = 9'o651;
		14'h83c: data = 9'o762;
		14'h83d: data = 9'o773;
		14'h83e: data = 9'o773;
		14'h83f: data = 9'o773;
		14'h840: data = 9'o773;
		14'h841: data = 9'o773;
		14'h842: data = 9'o773;
		14'h843: data = 9'o773;
		14'h844: data = 9'o773;
		14'h845: data = 9'o773;
		14'h846: data = 9'o773;
		14'h847: data = 9'o773;
		14'h848: data = 9'o773;
		14'h849: data = 9'o773;
		14'h84a: data = 9'o773;
		14'h84b: data = 9'o773;
		14'h84c: data = 9'o773;
		14'h84d: data = 9'o773;
		14'h84e: data = 9'o773;
		14'h84f: data = 9'o773;
		14'h850: data = 9'o773;
		14'h851: data = 9'o773;
		14'h852: data = 9'o773;
		14'h853: data = 9'o773;
		14'h854: data = 9'o773;
		14'h855: data = 9'o773;
		14'h856: data = 9'o773;
		14'h857: data = 9'o773;
		14'h858: data = 9'o773;
		14'h859: data = 9'o773;
		14'h85a: data = 9'o773;
		14'h85b: data = 9'o773;
		14'h85c: data = 9'o773;
		14'h85d: data = 9'o773;
		14'h85e: data = 9'o773;
		14'h85f: data = 9'o773;
		14'h860: data = 9'o773;
		14'h861: data = 9'o773;
		14'h862: data = 9'o773;
		14'h863: data = 9'o773;
		14'h864: data = 9'o252;
		14'h865: data = 9'o252;
		14'h866: data = 9'o773;
		14'h867: data = 9'o773;
		14'h868: data = 9'o773;
		14'h869: data = 9'o773;
		14'h86a: data = 9'o773;
		14'h86b: data = 9'o773;
		14'h86c: data = 9'o773;
		14'h86d: data = 9'o773;
		14'h86e: data = 9'o773;
		14'h86f: data = 9'o773;
		14'h870: data = 9'o773;
		14'h871: data = 9'o773;
		14'h872: data = 9'o773;
		14'h873: data = 9'o773;
		14'h874: data = 9'o773;
		14'h875: data = 9'o773;
		14'h876: data = 9'o773;
		14'h877: data = 9'o773;
		14'h878: data = 9'o773;
		14'h879: data = 9'o773;
		14'h87a: data = 9'o773;
		14'h87b: data = 9'o773;
		14'h87c: data = 9'o773;
		14'h87d: data = 9'o773;
		14'h87e: data = 9'o773;
		14'h87f: data = 9'o773;
		14'h880: data = 9'o773;
		14'h881: data = 9'o773;
		14'h882: data = 9'o773;
		14'h883: data = 9'o773;
		14'h884: data = 9'o773;
		14'h885: data = 9'o773;
		14'h886: data = 9'o773;
		14'h887: data = 9'o773;
		14'h888: data = 9'o773;
		14'h889: data = 9'o773;
		14'h88a: data = 9'o773;
		14'h88b: data = 9'o773;
		14'h88c: data = 9'o773;
		14'h88d: data = 9'o763;
		14'h88e: data = 9'o0;
		14'h88f: data = 9'o0;
		14'h890: data = 9'o0;
		14'h891: data = 9'o0;
		14'h892: data = 9'o0;
		14'h893: data = 9'o0;
		14'h894: data = 9'o0;
		14'h895: data = 9'o0;
		14'h896: data = 9'o0;
		14'h897: data = 9'o0;
		14'h898: data = 9'o0;
		14'h899: data = 9'o0;
		14'h89a: data = 9'o0;
		14'h89b: data = 9'o0;
		14'h89c: data = 9'o0;
		14'h89d: data = 9'o0;
		14'h89e: data = 9'o0;
		14'h89f: data = 9'o651;
		14'h8a0: data = 9'o762;
		14'h8a1: data = 9'o773;
		14'h8a2: data = 9'o773;
		14'h8a3: data = 9'o773;
		14'h8a4: data = 9'o773;
		14'h8a5: data = 9'o773;
		14'h8a6: data = 9'o773;
		14'h8a7: data = 9'o773;
		14'h8a8: data = 9'o773;
		14'h8a9: data = 9'o773;
		14'h8aa: data = 9'o773;
		14'h8ab: data = 9'o773;
		14'h8ac: data = 9'o773;
		14'h8ad: data = 9'o773;
		14'h8ae: data = 9'o773;
		14'h8af: data = 9'o773;
		14'h8b0: data = 9'o773;
		14'h8b1: data = 9'o773;
		14'h8b2: data = 9'o773;
		14'h8b3: data = 9'o773;
		14'h8b4: data = 9'o773;
		14'h8b5: data = 9'o773;
		14'h8b6: data = 9'o773;
		14'h8b7: data = 9'o773;
		14'h8b8: data = 9'o773;
		14'h8b9: data = 9'o773;
		14'h8ba: data = 9'o773;
		14'h8bb: data = 9'o773;
		14'h8bc: data = 9'o773;
		14'h8bd: data = 9'o773;
		14'h8be: data = 9'o773;
		14'h8bf: data = 9'o773;
		14'h8c0: data = 9'o773;
		14'h8c1: data = 9'o773;
		14'h8c2: data = 9'o773;
		14'h8c3: data = 9'o773;
		14'h8c4: data = 9'o773;
		14'h8c5: data = 9'o773;
		14'h8c6: data = 9'o773;
		14'h8c7: data = 9'o773;
		14'h8c8: data = 9'o252;
		14'h8c9: data = 9'o252;
		14'h8ca: data = 9'o673;
		14'h8cb: data = 9'o773;
		14'h8cc: data = 9'o773;
		14'h8cd: data = 9'o773;
		14'h8ce: data = 9'o773;
		14'h8cf: data = 9'o773;
		14'h8d0: data = 9'o773;
		14'h8d1: data = 9'o773;
		14'h8d2: data = 9'o773;
		14'h8d3: data = 9'o773;
		14'h8d4: data = 9'o773;
		14'h8d5: data = 9'o773;
		14'h8d6: data = 9'o773;
		14'h8d7: data = 9'o773;
		14'h8d8: data = 9'o773;
		14'h8d9: data = 9'o773;
		14'h8da: data = 9'o773;
		14'h8db: data = 9'o773;
		14'h8dc: data = 9'o773;
		14'h8dd: data = 9'o773;
		14'h8de: data = 9'o773;
		14'h8df: data = 9'o773;
		14'h8e0: data = 9'o773;
		14'h8e1: data = 9'o773;
		14'h8e2: data = 9'o773;
		14'h8e3: data = 9'o773;
		14'h8e4: data = 9'o773;
		14'h8e5: data = 9'o773;
		14'h8e6: data = 9'o773;
		14'h8e7: data = 9'o773;
		14'h8e8: data = 9'o773;
		14'h8e9: data = 9'o773;
		14'h8ea: data = 9'o773;
		14'h8eb: data = 9'o773;
		14'h8ec: data = 9'o773;
		14'h8ed: data = 9'o773;
		14'h8ee: data = 9'o773;
		14'h8ef: data = 9'o773;
		14'h8f0: data = 9'o773;
		14'h8f1: data = 9'o763;
		14'h8f2: data = 9'o0;
		14'h8f3: data = 9'o0;
		14'h8f4: data = 9'o0;
		14'h8f5: data = 9'o0;
		14'h8f6: data = 9'o0;
		14'h8f7: data = 9'o0;
		14'h8f8: data = 9'o0;
		14'h8f9: data = 9'o0;
		14'h8fa: data = 9'o0;
		14'h8fb: data = 9'o0;
		14'h8fc: data = 9'o0;
		14'h8fd: data = 9'o0;
		14'h8fe: data = 9'o0;
		14'h8ff: data = 9'o0;
		14'h900: data = 9'o0;
		14'h901: data = 9'o0;
		14'h902: data = 9'o0;
		14'h903: data = 9'o651;
		14'h904: data = 9'o762;
		14'h905: data = 9'o773;
		14'h906: data = 9'o773;
		14'h907: data = 9'o773;
		14'h908: data = 9'o773;
		14'h909: data = 9'o773;
		14'h90a: data = 9'o773;
		14'h90b: data = 9'o773;
		14'h90c: data = 9'o773;
		14'h90d: data = 9'o773;
		14'h90e: data = 9'o773;
		14'h90f: data = 9'o773;
		14'h910: data = 9'o773;
		14'h911: data = 9'o773;
		14'h912: data = 9'o773;
		14'h913: data = 9'o773;
		14'h914: data = 9'o773;
		14'h915: data = 9'o773;
		14'h916: data = 9'o773;
		14'h917: data = 9'o773;
		14'h918: data = 9'o773;
		14'h919: data = 9'o773;
		14'h91a: data = 9'o773;
		14'h91b: data = 9'o773;
		14'h91c: data = 9'o773;
		14'h91d: data = 9'o773;
		14'h91e: data = 9'o773;
		14'h91f: data = 9'o773;
		14'h920: data = 9'o773;
		14'h921: data = 9'o773;
		14'h922: data = 9'o773;
		14'h923: data = 9'o773;
		14'h924: data = 9'o773;
		14'h925: data = 9'o773;
		14'h926: data = 9'o773;
		14'h927: data = 9'o773;
		14'h928: data = 9'o773;
		14'h929: data = 9'o773;
		14'h92a: data = 9'o773;
		14'h92b: data = 9'o673;
		14'h92c: data = 9'o152;
		14'h92d: data = 9'o152;
		14'h92e: data = 9'o573;
		14'h92f: data = 9'o773;
		14'h930: data = 9'o773;
		14'h931: data = 9'o773;
		14'h932: data = 9'o773;
		14'h933: data = 9'o773;
		14'h934: data = 9'o773;
		14'h935: data = 9'o773;
		14'h936: data = 9'o773;
		14'h937: data = 9'o773;
		14'h938: data = 9'o773;
		14'h939: data = 9'o773;
		14'h93a: data = 9'o773;
		14'h93b: data = 9'o773;
		14'h93c: data = 9'o773;
		14'h93d: data = 9'o773;
		14'h93e: data = 9'o773;
		14'h93f: data = 9'o773;
		14'h940: data = 9'o773;
		14'h941: data = 9'o773;
		14'h942: data = 9'o773;
		14'h943: data = 9'o773;
		14'h944: data = 9'o773;
		14'h945: data = 9'o773;
		14'h946: data = 9'o773;
		14'h947: data = 9'o773;
		14'h948: data = 9'o773;
		14'h949: data = 9'o773;
		14'h94a: data = 9'o773;
		14'h94b: data = 9'o773;
		14'h94c: data = 9'o773;
		14'h94d: data = 9'o773;
		14'h94e: data = 9'o773;
		14'h94f: data = 9'o773;
		14'h950: data = 9'o773;
		14'h951: data = 9'o773;
		14'h952: data = 9'o773;
		14'h953: data = 9'o773;
		14'h954: data = 9'o773;
		14'h955: data = 9'o763;
		14'h956: data = 9'o0;
		14'h957: data = 9'o0;
		14'h958: data = 9'o0;
		14'h959: data = 9'o0;
		14'h95a: data = 9'o0;
		14'h95b: data = 9'o0;
		14'h95c: data = 9'o0;
		14'h95d: data = 9'o0;
		14'h95e: data = 9'o0;
		14'h95f: data = 9'o0;
		14'h960: data = 9'o0;
		14'h961: data = 9'o0;
		14'h962: data = 9'o0;
		14'h963: data = 9'o0;
		14'h964: data = 9'o0;
		14'h965: data = 9'o0;
		14'h966: data = 9'o0;
		14'h967: data = 9'o551;
		14'h968: data = 9'o762;
		14'h969: data = 9'o773;
		14'h96a: data = 9'o773;
		14'h96b: data = 9'o773;
		14'h96c: data = 9'o773;
		14'h96d: data = 9'o773;
		14'h96e: data = 9'o773;
		14'h96f: data = 9'o773;
		14'h970: data = 9'o773;
		14'h971: data = 9'o773;
		14'h972: data = 9'o773;
		14'h973: data = 9'o773;
		14'h974: data = 9'o773;
		14'h975: data = 9'o773;
		14'h976: data = 9'o773;
		14'h977: data = 9'o773;
		14'h978: data = 9'o773;
		14'h979: data = 9'o773;
		14'h97a: data = 9'o773;
		14'h97b: data = 9'o773;
		14'h97c: data = 9'o773;
		14'h97d: data = 9'o773;
		14'h97e: data = 9'o773;
		14'h97f: data = 9'o773;
		14'h980: data = 9'o773;
		14'h981: data = 9'o773;
		14'h982: data = 9'o773;
		14'h983: data = 9'o773;
		14'h984: data = 9'o773;
		14'h985: data = 9'o773;
		14'h986: data = 9'o773;
		14'h987: data = 9'o773;
		14'h988: data = 9'o773;
		14'h989: data = 9'o773;
		14'h98a: data = 9'o773;
		14'h98b: data = 9'o773;
		14'h98c: data = 9'o773;
		14'h98d: data = 9'o773;
		14'h98e: data = 9'o773;
		14'h98f: data = 9'o463;
		14'h990: data = 9'o152;
		14'h991: data = 9'o152;
		14'h992: data = 9'o463;
		14'h993: data = 9'o773;
		14'h994: data = 9'o773;
		14'h995: data = 9'o773;
		14'h996: data = 9'o773;
		14'h997: data = 9'o773;
		14'h998: data = 9'o773;
		14'h999: data = 9'o773;
		14'h99a: data = 9'o773;
		14'h99b: data = 9'o773;
		14'h99c: data = 9'o773;
		14'h99d: data = 9'o773;
		14'h99e: data = 9'o773;
		14'h99f: data = 9'o773;
		14'h9a0: data = 9'o773;
		14'h9a1: data = 9'o773;
		14'h9a2: data = 9'o773;
		14'h9a3: data = 9'o773;
		14'h9a4: data = 9'o773;
		14'h9a5: data = 9'o773;
		14'h9a6: data = 9'o773;
		14'h9a7: data = 9'o773;
		14'h9a8: data = 9'o773;
		14'h9a9: data = 9'o773;
		14'h9aa: data = 9'o773;
		14'h9ab: data = 9'o773;
		14'h9ac: data = 9'o773;
		14'h9ad: data = 9'o773;
		14'h9ae: data = 9'o773;
		14'h9af: data = 9'o773;
		14'h9b0: data = 9'o773;
		14'h9b1: data = 9'o773;
		14'h9b2: data = 9'o773;
		14'h9b3: data = 9'o773;
		14'h9b4: data = 9'o773;
		14'h9b5: data = 9'o773;
		14'h9b6: data = 9'o773;
		14'h9b7: data = 9'o773;
		14'h9b8: data = 9'o773;
		14'h9b9: data = 9'o763;
		14'h9ba: data = 9'o0;
		14'h9bb: data = 9'o0;
		14'h9bc: data = 9'o0;
		14'h9bd: data = 9'o0;
		14'h9be: data = 9'o0;
		14'h9bf: data = 9'o0;
		14'h9c0: data = 9'o0;
		14'h9c1: data = 9'o0;
		14'h9c2: data = 9'o0;
		14'h9c3: data = 9'o0;
		14'h9c4: data = 9'o0;
		14'h9c5: data = 9'o0;
		14'h9c6: data = 9'o0;
		14'h9c7: data = 9'o0;
		14'h9c8: data = 9'o0;
		14'h9c9: data = 9'o0;
		14'h9ca: data = 9'o0;
		14'h9cb: data = 9'o551;
		14'h9cc: data = 9'o762;
		14'h9cd: data = 9'o773;
		14'h9ce: data = 9'o773;
		14'h9cf: data = 9'o773;
		14'h9d0: data = 9'o773;
		14'h9d1: data = 9'o773;
		14'h9d2: data = 9'o773;
		14'h9d3: data = 9'o773;
		14'h9d4: data = 9'o773;
		14'h9d5: data = 9'o773;
		14'h9d6: data = 9'o773;
		14'h9d7: data = 9'o773;
		14'h9d8: data = 9'o773;
		14'h9d9: data = 9'o773;
		14'h9da: data = 9'o773;
		14'h9db: data = 9'o773;
		14'h9dc: data = 9'o773;
		14'h9dd: data = 9'o773;
		14'h9de: data = 9'o773;
		14'h9df: data = 9'o773;
		14'h9e0: data = 9'o773;
		14'h9e1: data = 9'o773;
		14'h9e2: data = 9'o773;
		14'h9e3: data = 9'o773;
		14'h9e4: data = 9'o773;
		14'h9e5: data = 9'o773;
		14'h9e6: data = 9'o773;
		14'h9e7: data = 9'o773;
		14'h9e8: data = 9'o773;
		14'h9e9: data = 9'o773;
		14'h9ea: data = 9'o773;
		14'h9eb: data = 9'o773;
		14'h9ec: data = 9'o773;
		14'h9ed: data = 9'o773;
		14'h9ee: data = 9'o773;
		14'h9ef: data = 9'o773;
		14'h9f0: data = 9'o773;
		14'h9f1: data = 9'o773;
		14'h9f2: data = 9'o773;
		14'h9f3: data = 9'o352;
		14'h9f4: data = 9'o152;
		14'h9f5: data = 9'o152;
		14'h9f6: data = 9'o252;
		14'h9f7: data = 9'o673;
		14'h9f8: data = 9'o773;
		14'h9f9: data = 9'o773;
		14'h9fa: data = 9'o773;
		14'h9fb: data = 9'o773;
		14'h9fc: data = 9'o773;
		14'h9fd: data = 9'o773;
		14'h9fe: data = 9'o773;
		14'h9ff: data = 9'o773;
		14'ha00: data = 9'o773;
		14'ha01: data = 9'o773;
		14'ha02: data = 9'o773;
		14'ha03: data = 9'o773;
		14'ha04: data = 9'o773;
		14'ha05: data = 9'o773;
		14'ha06: data = 9'o773;
		14'ha07: data = 9'o773;
		14'ha08: data = 9'o773;
		14'ha09: data = 9'o773;
		14'ha0a: data = 9'o773;
		14'ha0b: data = 9'o773;
		14'ha0c: data = 9'o773;
		14'ha0d: data = 9'o773;
		14'ha0e: data = 9'o773;
		14'ha0f: data = 9'o773;
		14'ha10: data = 9'o773;
		14'ha11: data = 9'o773;
		14'ha12: data = 9'o773;
		14'ha13: data = 9'o773;
		14'ha14: data = 9'o773;
		14'ha15: data = 9'o773;
		14'ha16: data = 9'o773;
		14'ha17: data = 9'o773;
		14'ha18: data = 9'o773;
		14'ha19: data = 9'o773;
		14'ha1a: data = 9'o773;
		14'ha1b: data = 9'o773;
		14'ha1c: data = 9'o773;
		14'ha1d: data = 9'o762;
		14'ha1e: data = 9'o0;
		14'ha1f: data = 9'o0;
		14'ha20: data = 9'o0;
		14'ha21: data = 9'o0;
		14'ha22: data = 9'o0;
		14'ha23: data = 9'o0;
		14'ha24: data = 9'o0;
		14'ha25: data = 9'o0;
		14'ha26: data = 9'o0;
		14'ha27: data = 9'o0;
		14'ha28: data = 9'o0;
		14'ha29: data = 9'o0;
		14'ha2a: data = 9'o0;
		14'ha2b: data = 9'o0;
		14'ha2c: data = 9'o0;
		14'ha2d: data = 9'o0;
		14'ha2e: data = 9'o0;
		14'ha2f: data = 9'o551;
		14'ha30: data = 9'o762;
		14'ha31: data = 9'o773;
		14'ha32: data = 9'o773;
		14'ha33: data = 9'o773;
		14'ha34: data = 9'o773;
		14'ha35: data = 9'o773;
		14'ha36: data = 9'o773;
		14'ha37: data = 9'o773;
		14'ha38: data = 9'o773;
		14'ha39: data = 9'o773;
		14'ha3a: data = 9'o773;
		14'ha3b: data = 9'o773;
		14'ha3c: data = 9'o773;
		14'ha3d: data = 9'o773;
		14'ha3e: data = 9'o773;
		14'ha3f: data = 9'o773;
		14'ha40: data = 9'o773;
		14'ha41: data = 9'o773;
		14'ha42: data = 9'o773;
		14'ha43: data = 9'o773;
		14'ha44: data = 9'o773;
		14'ha45: data = 9'o773;
		14'ha46: data = 9'o773;
		14'ha47: data = 9'o773;
		14'ha48: data = 9'o773;
		14'ha49: data = 9'o773;
		14'ha4a: data = 9'o773;
		14'ha4b: data = 9'o773;
		14'ha4c: data = 9'o773;
		14'ha4d: data = 9'o773;
		14'ha4e: data = 9'o773;
		14'ha4f: data = 9'o773;
		14'ha50: data = 9'o773;
		14'ha51: data = 9'o773;
		14'ha52: data = 9'o773;
		14'ha53: data = 9'o773;
		14'ha54: data = 9'o773;
		14'ha55: data = 9'o773;
		14'ha56: data = 9'o673;
		14'ha57: data = 9'o252;
		14'ha58: data = 9'o152;
		14'ha59: data = 9'o152;
		14'ha5a: data = 9'o252;
		14'ha5b: data = 9'o673;
		14'ha5c: data = 9'o773;
		14'ha5d: data = 9'o773;
		14'ha5e: data = 9'o773;
		14'ha5f: data = 9'o773;
		14'ha60: data = 9'o773;
		14'ha61: data = 9'o773;
		14'ha62: data = 9'o773;
		14'ha63: data = 9'o773;
		14'ha64: data = 9'o773;
		14'ha65: data = 9'o773;
		14'ha66: data = 9'o773;
		14'ha67: data = 9'o773;
		14'ha68: data = 9'o773;
		14'ha69: data = 9'o773;
		14'ha6a: data = 9'o773;
		14'ha6b: data = 9'o773;
		14'ha6c: data = 9'o773;
		14'ha6d: data = 9'o773;
		14'ha6e: data = 9'o773;
		14'ha6f: data = 9'o773;
		14'ha70: data = 9'o773;
		14'ha71: data = 9'o773;
		14'ha72: data = 9'o773;
		14'ha73: data = 9'o773;
		14'ha74: data = 9'o773;
		14'ha75: data = 9'o773;
		14'ha76: data = 9'o773;
		14'ha77: data = 9'o773;
		14'ha78: data = 9'o773;
		14'ha79: data = 9'o773;
		14'ha7a: data = 9'o773;
		14'ha7b: data = 9'o773;
		14'ha7c: data = 9'o773;
		14'ha7d: data = 9'o773;
		14'ha7e: data = 9'o773;
		14'ha7f: data = 9'o773;
		14'ha80: data = 9'o773;
		14'ha81: data = 9'o762;
		14'ha82: data = 9'o0;
		14'ha83: data = 9'o0;
		14'ha84: data = 9'o0;
		14'ha85: data = 9'o0;
		14'ha86: data = 9'o0;
		14'ha87: data = 9'o0;
		14'ha88: data = 9'o0;
		14'ha89: data = 9'o0;
		14'ha8a: data = 9'o0;
		14'ha8b: data = 9'o0;
		14'ha8c: data = 9'o0;
		14'ha8d: data = 9'o0;
		14'ha8e: data = 9'o0;
		14'ha8f: data = 9'o0;
		14'ha90: data = 9'o0;
		14'ha91: data = 9'o0;
		14'ha92: data = 9'o0;
		14'ha93: data = 9'o651;
		14'ha94: data = 9'o762;
		14'ha95: data = 9'o773;
		14'ha96: data = 9'o773;
		14'ha97: data = 9'o773;
		14'ha98: data = 9'o773;
		14'ha99: data = 9'o773;
		14'ha9a: data = 9'o773;
		14'ha9b: data = 9'o773;
		14'ha9c: data = 9'o773;
		14'ha9d: data = 9'o773;
		14'ha9e: data = 9'o773;
		14'ha9f: data = 9'o773;
		14'haa0: data = 9'o773;
		14'haa1: data = 9'o773;
		14'haa2: data = 9'o773;
		14'haa3: data = 9'o773;
		14'haa4: data = 9'o773;
		14'haa5: data = 9'o773;
		14'haa6: data = 9'o773;
		14'haa7: data = 9'o773;
		14'haa8: data = 9'o773;
		14'haa9: data = 9'o773;
		14'haaa: data = 9'o773;
		14'haab: data = 9'o773;
		14'haac: data = 9'o773;
		14'haad: data = 9'o773;
		14'haae: data = 9'o773;
		14'haaf: data = 9'o773;
		14'hab0: data = 9'o773;
		14'hab1: data = 9'o773;
		14'hab2: data = 9'o773;
		14'hab3: data = 9'o773;
		14'hab4: data = 9'o773;
		14'hab5: data = 9'o773;
		14'hab6: data = 9'o773;
		14'hab7: data = 9'o773;
		14'hab8: data = 9'o773;
		14'hab9: data = 9'o773;
		14'haba: data = 9'o573;
		14'habb: data = 9'o252;
		14'habc: data = 9'o152;
		14'habd: data = 9'o152;
		14'habe: data = 9'o252;
		14'habf: data = 9'o573;
		14'hac0: data = 9'o773;
		14'hac1: data = 9'o773;
		14'hac2: data = 9'o773;
		14'hac3: data = 9'o773;
		14'hac4: data = 9'o773;
		14'hac5: data = 9'o773;
		14'hac6: data = 9'o773;
		14'hac7: data = 9'o773;
		14'hac8: data = 9'o773;
		14'hac9: data = 9'o773;
		14'haca: data = 9'o773;
		14'hacb: data = 9'o773;
		14'hacc: data = 9'o773;
		14'hacd: data = 9'o773;
		14'hace: data = 9'o773;
		14'hacf: data = 9'o773;
		14'had0: data = 9'o773;
		14'had1: data = 9'o773;
		14'had2: data = 9'o773;
		14'had3: data = 9'o773;
		14'had4: data = 9'o773;
		14'had5: data = 9'o773;
		14'had6: data = 9'o773;
		14'had7: data = 9'o773;
		14'had8: data = 9'o773;
		14'had9: data = 9'o773;
		14'hada: data = 9'o773;
		14'hadb: data = 9'o773;
		14'hadc: data = 9'o773;
		14'hadd: data = 9'o773;
		14'hade: data = 9'o773;
		14'hadf: data = 9'o773;
		14'hae0: data = 9'o773;
		14'hae1: data = 9'o773;
		14'hae2: data = 9'o773;
		14'hae3: data = 9'o773;
		14'hae4: data = 9'o773;
		14'hae5: data = 9'o762;
		14'hae6: data = 9'o0;
		14'hae7: data = 9'o0;
		14'hae8: data = 9'o0;
		14'hae9: data = 9'o0;
		14'haea: data = 9'o0;
		14'haeb: data = 9'o0;
		14'haec: data = 9'o0;
		14'haed: data = 9'o0;
		14'haee: data = 9'o0;
		14'haef: data = 9'o0;
		14'haf0: data = 9'o0;
		14'haf1: data = 9'o0;
		14'haf2: data = 9'o0;
		14'haf3: data = 9'o0;
		14'haf4: data = 9'o0;
		14'haf5: data = 9'o0;
		14'haf6: data = 9'o0;
		14'haf7: data = 9'o641;
		14'haf8: data = 9'o762;
		14'haf9: data = 9'o773;
		14'hafa: data = 9'o773;
		14'hafb: data = 9'o673;
		14'hafc: data = 9'o773;
		14'hafd: data = 9'o773;
		14'hafe: data = 9'o773;
		14'haff: data = 9'o773;
		14'hb00: data = 9'o773;
		14'hb01: data = 9'o773;
		14'hb02: data = 9'o673;
		14'hb03: data = 9'o773;
		14'hb04: data = 9'o773;
		14'hb05: data = 9'o773;
		14'hb06: data = 9'o773;
		14'hb07: data = 9'o773;
		14'hb08: data = 9'o773;
		14'hb09: data = 9'o773;
		14'hb0a: data = 9'o773;
		14'hb0b: data = 9'o773;
		14'hb0c: data = 9'o773;
		14'hb0d: data = 9'o773;
		14'hb0e: data = 9'o773;
		14'hb0f: data = 9'o773;
		14'hb10: data = 9'o773;
		14'hb11: data = 9'o773;
		14'hb12: data = 9'o773;
		14'hb13: data = 9'o773;
		14'hb14: data = 9'o773;
		14'hb15: data = 9'o773;
		14'hb16: data = 9'o773;
		14'hb17: data = 9'o773;
		14'hb18: data = 9'o773;
		14'hb19: data = 9'o773;
		14'hb1a: data = 9'o773;
		14'hb1b: data = 9'o773;
		14'hb1c: data = 9'o773;
		14'hb1d: data = 9'o773;
		14'hb1e: data = 9'o473;
		14'hb1f: data = 9'o142;
		14'hb20: data = 9'o152;
		14'hb21: data = 9'o152;
		14'hb22: data = 9'o142;
		14'hb23: data = 9'o463;
		14'hb24: data = 9'o773;
		14'hb25: data = 9'o773;
		14'hb26: data = 9'o773;
		14'hb27: data = 9'o773;
		14'hb28: data = 9'o773;
		14'hb29: data = 9'o773;
		14'hb2a: data = 9'o773;
		14'hb2b: data = 9'o773;
		14'hb2c: data = 9'o773;
		14'hb2d: data = 9'o773;
		14'hb2e: data = 9'o773;
		14'hb2f: data = 9'o773;
		14'hb30: data = 9'o773;
		14'hb31: data = 9'o773;
		14'hb32: data = 9'o773;
		14'hb33: data = 9'o773;
		14'hb34: data = 9'o773;
		14'hb35: data = 9'o773;
		14'hb36: data = 9'o773;
		14'hb37: data = 9'o773;
		14'hb38: data = 9'o773;
		14'hb39: data = 9'o773;
		14'hb3a: data = 9'o773;
		14'hb3b: data = 9'o773;
		14'hb3c: data = 9'o773;
		14'hb3d: data = 9'o773;
		14'hb3e: data = 9'o773;
		14'hb3f: data = 9'o773;
		14'hb40: data = 9'o773;
		14'hb41: data = 9'o773;
		14'hb42: data = 9'o773;
		14'hb43: data = 9'o773;
		14'hb44: data = 9'o773;
		14'hb45: data = 9'o773;
		14'hb46: data = 9'o673;
		14'hb47: data = 9'o673;
		14'hb48: data = 9'o773;
		14'hb49: data = 9'o762;
		14'hb4a: data = 9'o0;
		14'hb4b: data = 9'o0;
		14'hb4c: data = 9'o0;
		14'hb4d: data = 9'o0;
		14'hb4e: data = 9'o0;
		14'hb4f: data = 9'o0;
		14'hb50: data = 9'o0;
		14'hb51: data = 9'o0;
		14'hb52: data = 9'o0;
		14'hb53: data = 9'o0;
		14'hb54: data = 9'o0;
		14'hb55: data = 9'o0;
		14'hb56: data = 9'o0;
		14'hb57: data = 9'o0;
		14'hb58: data = 9'o0;
		14'hb59: data = 9'o0;
		14'hb5a: data = 9'o0;
		14'hb5b: data = 9'o651;
		14'hb5c: data = 9'o762;
		14'hb5d: data = 9'o773;
		14'hb5e: data = 9'o352;
		14'hb5f: data = 9'o252;
		14'hb60: data = 9'o252;
		14'hb61: data = 9'o362;
		14'hb62: data = 9'o773;
		14'hb63: data = 9'o773;
		14'hb64: data = 9'o673;
		14'hb65: data = 9'o352;
		14'hb66: data = 9'o252;
		14'hb67: data = 9'o352;
		14'hb68: data = 9'o673;
		14'hb69: data = 9'o773;
		14'hb6a: data = 9'o773;
		14'hb6b: data = 9'o563;
		14'hb6c: data = 9'o252;
		14'hb6d: data = 9'o252;
		14'hb6e: data = 9'o563;
		14'hb6f: data = 9'o773;
		14'hb70: data = 9'o773;
		14'hb71: data = 9'o673;
		14'hb72: data = 9'o252;
		14'hb73: data = 9'o252;
		14'hb74: data = 9'o252;
		14'hb75: data = 9'o352;
		14'hb76: data = 9'o673;
		14'hb77: data = 9'o773;
		14'hb78: data = 9'o773;
		14'hb79: data = 9'o773;
		14'hb7a: data = 9'o773;
		14'hb7b: data = 9'o773;
		14'hb7c: data = 9'o773;
		14'hb7d: data = 9'o773;
		14'hb7e: data = 9'o773;
		14'hb7f: data = 9'o773;
		14'hb80: data = 9'o773;
		14'hb81: data = 9'o773;
		14'hb82: data = 9'o363;
		14'hb83: data = 9'o152;
		14'hb84: data = 9'o152;
		14'hb85: data = 9'o152;
		14'hb86: data = 9'o142;
		14'hb87: data = 9'o353;
		14'hb88: data = 9'o773;
		14'hb89: data = 9'o773;
		14'hb8a: data = 9'o773;
		14'hb8b: data = 9'o773;
		14'hb8c: data = 9'o773;
		14'hb8d: data = 9'o773;
		14'hb8e: data = 9'o773;
		14'hb8f: data = 9'o773;
		14'hb90: data = 9'o773;
		14'hb91: data = 9'o773;
		14'hb92: data = 9'o773;
		14'hb93: data = 9'o673;
		14'hb94: data = 9'o252;
		14'hb95: data = 9'o252;
		14'hb96: data = 9'o252;
		14'hb97: data = 9'o252;
		14'hb98: data = 9'o673;
		14'hb99: data = 9'o773;
		14'hb9a: data = 9'o773;
		14'hb9b: data = 9'o573;
		14'hb9c: data = 9'o252;
		14'hb9d: data = 9'o252;
		14'hb9e: data = 9'o463;
		14'hb9f: data = 9'o773;
		14'hba0: data = 9'o773;
		14'hba1: data = 9'o673;
		14'hba2: data = 9'o352;
		14'hba3: data = 9'o252;
		14'hba4: data = 9'o352;
		14'hba5: data = 9'o773;
		14'hba6: data = 9'o773;
		14'hba7: data = 9'o773;
		14'hba8: data = 9'o463;
		14'hba9: data = 9'o252;
		14'hbaa: data = 9'o252;
		14'hbab: data = 9'o352;
		14'hbac: data = 9'o773;
		14'hbad: data = 9'o662;
		14'hbae: data = 9'o0;
		14'hbaf: data = 9'o0;
		14'hbb0: data = 9'o0;
		14'hbb1: data = 9'o0;
		14'hbb2: data = 9'o0;
		14'hbb3: data = 9'o0;
		14'hbb4: data = 9'o0;
		14'hbb5: data = 9'o0;
		14'hbb6: data = 9'o0;
		14'hbb7: data = 9'o0;
		14'hbb8: data = 9'o0;
		14'hbb9: data = 9'o0;
		14'hbba: data = 9'o0;
		14'hbbb: data = 9'o0;
		14'hbbc: data = 9'o0;
		14'hbbd: data = 9'o0;
		14'hbbe: data = 9'o0;
		14'hbbf: data = 9'o551;
		14'hbc0: data = 9'o762;
		14'hbc1: data = 9'o773;
		14'hbc2: data = 9'o252;
		14'hbc3: data = 9'o152;
		14'hbc4: data = 9'o152;
		14'hbc5: data = 9'o363;
		14'hbc6: data = 9'o673;
		14'hbc7: data = 9'o773;
		14'hbc8: data = 9'o773;
		14'hbc9: data = 9'o352;
		14'hbca: data = 9'o152;
		14'hbcb: data = 9'o252;
		14'hbcc: data = 9'o673;
		14'hbcd: data = 9'o773;
		14'hbce: data = 9'o773;
		14'hbcf: data = 9'o463;
		14'hbd0: data = 9'o152;
		14'hbd1: data = 9'o152;
		14'hbd2: data = 9'o463;
		14'hbd3: data = 9'o773;
		14'hbd4: data = 9'o773;
		14'hbd5: data = 9'o673;
		14'hbd6: data = 9'o152;
		14'hbd7: data = 9'o152;
		14'hbd8: data = 9'o152;
		14'hbd9: data = 9'o252;
		14'hbda: data = 9'o573;
		14'hbdb: data = 9'o773;
		14'hbdc: data = 9'o773;
		14'hbdd: data = 9'o773;
		14'hbde: data = 9'o773;
		14'hbdf: data = 9'o773;
		14'hbe0: data = 9'o773;
		14'hbe1: data = 9'o773;
		14'hbe2: data = 9'o773;
		14'hbe3: data = 9'o773;
		14'hbe4: data = 9'o773;
		14'hbe5: data = 9'o673;
		14'hbe6: data = 9'o252;
		14'hbe7: data = 9'o152;
		14'hbe8: data = 9'o152;
		14'hbe9: data = 9'o152;
		14'hbea: data = 9'o152;
		14'hbeb: data = 9'o252;
		14'hbec: data = 9'o673;
		14'hbed: data = 9'o773;
		14'hbee: data = 9'o773;
		14'hbef: data = 9'o773;
		14'hbf0: data = 9'o773;
		14'hbf1: data = 9'o773;
		14'hbf2: data = 9'o773;
		14'hbf3: data = 9'o773;
		14'hbf4: data = 9'o773;
		14'hbf5: data = 9'o773;
		14'hbf6: data = 9'o773;
		14'hbf7: data = 9'o673;
		14'hbf8: data = 9'o152;
		14'hbf9: data = 9'o152;
		14'hbfa: data = 9'o152;
		14'hbfb: data = 9'o142;
		14'hbfc: data = 9'o673;
		14'hbfd: data = 9'o773;
		14'hbfe: data = 9'o673;
		14'hbff: data = 9'o463;
		14'hc00: data = 9'o152;
		14'hc01: data = 9'o152;
		14'hc02: data = 9'o463;
		14'hc03: data = 9'o673;
		14'hc04: data = 9'o773;
		14'hc05: data = 9'o673;
		14'hc06: data = 9'o252;
		14'hc07: data = 9'o142;
		14'hc08: data = 9'o252;
		14'hc09: data = 9'o673;
		14'hc0a: data = 9'o773;
		14'hc0b: data = 9'o773;
		14'hc0c: data = 9'o362;
		14'hc0d: data = 9'o152;
		14'hc0e: data = 9'o152;
		14'hc0f: data = 9'o252;
		14'hc10: data = 9'o773;
		14'hc11: data = 9'o763;
		14'hc12: data = 9'o0;
		14'hc13: data = 9'o0;
		14'hc14: data = 9'o0;
		14'hc15: data = 9'o0;
		14'hc16: data = 9'o0;
		14'hc17: data = 9'o0;
		14'hc18: data = 9'o0;
		14'hc19: data = 9'o0;
		14'hc1a: data = 9'o0;
		14'hc1b: data = 9'o0;
		14'hc1c: data = 9'o0;
		14'hc1d: data = 9'o0;
		14'hc1e: data = 9'o0;
		14'hc1f: data = 9'o0;
		14'hc20: data = 9'o0;
		14'hc21: data = 9'o0;
		14'hc22: data = 9'o0;
		14'hc23: data = 9'o651;
		14'hc24: data = 9'o762;
		14'hc25: data = 9'o773;
		14'hc26: data = 9'o252;
		14'hc27: data = 9'o152;
		14'hc28: data = 9'o152;
		14'hc29: data = 9'o263;
		14'hc2a: data = 9'o673;
		14'hc2b: data = 9'o773;
		14'hc2c: data = 9'o773;
		14'hc2d: data = 9'o352;
		14'hc2e: data = 9'o152;
		14'hc2f: data = 9'o252;
		14'hc30: data = 9'o673;
		14'hc31: data = 9'o773;
		14'hc32: data = 9'o773;
		14'hc33: data = 9'o463;
		14'hc34: data = 9'o152;
		14'hc35: data = 9'o152;
		14'hc36: data = 9'o463;
		14'hc37: data = 9'o773;
		14'hc38: data = 9'o773;
		14'hc39: data = 9'o673;
		14'hc3a: data = 9'o152;
		14'hc3b: data = 9'o52;
		14'hc3c: data = 9'o152;
		14'hc3d: data = 9'o152;
		14'hc3e: data = 9'o573;
		14'hc3f: data = 9'o773;
		14'hc40: data = 9'o773;
		14'hc41: data = 9'o773;
		14'hc42: data = 9'o773;
		14'hc43: data = 9'o773;
		14'hc44: data = 9'o773;
		14'hc45: data = 9'o773;
		14'hc46: data = 9'o773;
		14'hc47: data = 9'o773;
		14'hc48: data = 9'o773;
		14'hc49: data = 9'o673;
		14'hc4a: data = 9'o252;
		14'hc4b: data = 9'o152;
		14'hc4c: data = 9'o152;
		14'hc4d: data = 9'o152;
		14'hc4e: data = 9'o152;
		14'hc4f: data = 9'o152;
		14'hc50: data = 9'o673;
		14'hc51: data = 9'o773;
		14'hc52: data = 9'o773;
		14'hc53: data = 9'o773;
		14'hc54: data = 9'o773;
		14'hc55: data = 9'o773;
		14'hc56: data = 9'o773;
		14'hc57: data = 9'o773;
		14'hc58: data = 9'o773;
		14'hc59: data = 9'o773;
		14'hc5a: data = 9'o773;
		14'hc5b: data = 9'o673;
		14'hc5c: data = 9'o142;
		14'hc5d: data = 9'o52;
		14'hc5e: data = 9'o152;
		14'hc5f: data = 9'o152;
		14'hc60: data = 9'o573;
		14'hc61: data = 9'o673;
		14'hc62: data = 9'o773;
		14'hc63: data = 9'o573;
		14'hc64: data = 9'o152;
		14'hc65: data = 9'o152;
		14'hc66: data = 9'o463;
		14'hc67: data = 9'o673;
		14'hc68: data = 9'o773;
		14'hc69: data = 9'o673;
		14'hc6a: data = 9'o252;
		14'hc6b: data = 9'o152;
		14'hc6c: data = 9'o352;
		14'hc6d: data = 9'o673;
		14'hc6e: data = 9'o773;
		14'hc6f: data = 9'o773;
		14'hc70: data = 9'o363;
		14'hc71: data = 9'o152;
		14'hc72: data = 9'o152;
		14'hc73: data = 9'o252;
		14'hc74: data = 9'o773;
		14'hc75: data = 9'o662;
		14'hc76: data = 9'o0;
		14'hc77: data = 9'o0;
		14'hc78: data = 9'o0;
		14'hc79: data = 9'o0;
		14'hc7a: data = 9'o0;
		14'hc7b: data = 9'o0;
		14'hc7c: data = 9'o0;
		14'hc7d: data = 9'o0;
		14'hc7e: data = 9'o0;
		14'hc7f: data = 9'o0;
		14'hc80: data = 9'o0;
		14'hc81: data = 9'o0;
		14'hc82: data = 9'o0;
		14'hc83: data = 9'o0;
		14'hc84: data = 9'o0;
		14'hc85: data = 9'o0;
		14'hc86: data = 9'o0;
		14'hc87: data = 9'o651;
		14'hc88: data = 9'o762;
		14'hc89: data = 9'o773;
		14'hc8a: data = 9'o252;
		14'hc8b: data = 9'o152;
		14'hc8c: data = 9'o52;
		14'hc8d: data = 9'o263;
		14'hc8e: data = 9'o573;
		14'hc8f: data = 9'o573;
		14'hc90: data = 9'o573;
		14'hc91: data = 9'o252;
		14'hc92: data = 9'o152;
		14'hc93: data = 9'o152;
		14'hc94: data = 9'o473;
		14'hc95: data = 9'o563;
		14'hc96: data = 9'o573;
		14'hc97: data = 9'o363;
		14'hc98: data = 9'o152;
		14'hc99: data = 9'o152;
		14'hc9a: data = 9'o363;
		14'hc9b: data = 9'o573;
		14'hc9c: data = 9'o573;
		14'hc9d: data = 9'o463;
		14'hc9e: data = 9'o152;
		14'hc9f: data = 9'o52;
		14'hca0: data = 9'o52;
		14'hca1: data = 9'o152;
		14'hca2: data = 9'o673;
		14'hca3: data = 9'o773;
		14'hca4: data = 9'o773;
		14'hca5: data = 9'o773;
		14'hca6: data = 9'o773;
		14'hca7: data = 9'o773;
		14'hca8: data = 9'o773;
		14'hca9: data = 9'o773;
		14'hcaa: data = 9'o773;
		14'hcab: data = 9'o773;
		14'hcac: data = 9'o773;
		14'hcad: data = 9'o573;
		14'hcae: data = 9'o152;
		14'hcaf: data = 9'o152;
		14'hcb0: data = 9'o152;
		14'hcb1: data = 9'o152;
		14'hcb2: data = 9'o152;
		14'hcb3: data = 9'o152;
		14'hcb4: data = 9'o573;
		14'hcb5: data = 9'o773;
		14'hcb6: data = 9'o773;
		14'hcb7: data = 9'o773;
		14'hcb8: data = 9'o773;
		14'hcb9: data = 9'o773;
		14'hcba: data = 9'o773;
		14'hcbb: data = 9'o773;
		14'hcbc: data = 9'o773;
		14'hcbd: data = 9'o773;
		14'hcbe: data = 9'o773;
		14'hcbf: data = 9'o673;
		14'hcc0: data = 9'o152;
		14'hcc1: data = 9'o52;
		14'hcc2: data = 9'o52;
		14'hcc3: data = 9'o152;
		14'hcc4: data = 9'o473;
		14'hcc5: data = 9'o573;
		14'hcc6: data = 9'o573;
		14'hcc7: data = 9'o463;
		14'hcc8: data = 9'o142;
		14'hcc9: data = 9'o152;
		14'hcca: data = 9'o353;
		14'hccb: data = 9'o573;
		14'hccc: data = 9'o573;
		14'hccd: data = 9'o473;
		14'hcce: data = 9'o152;
		14'hccf: data = 9'o142;
		14'hcd0: data = 9'o252;
		14'hcd1: data = 9'o573;
		14'hcd2: data = 9'o573;
		14'hcd3: data = 9'o573;
		14'hcd4: data = 9'o263;
		14'hcd5: data = 9'o52;
		14'hcd6: data = 9'o152;
		14'hcd7: data = 9'o252;
		14'hcd8: data = 9'o773;
		14'hcd9: data = 9'o762;
		14'hcda: data = 9'o0;
		14'hcdb: data = 9'o0;
		14'hcdc: data = 9'o0;
		14'hcdd: data = 9'o0;
		14'hcde: data = 9'o0;
		14'hcdf: data = 9'o0;
		14'hce0: data = 9'o0;
		14'hce1: data = 9'o0;
		14'hce2: data = 9'o0;
		14'hce3: data = 9'o0;
		14'hce4: data = 9'o0;
		14'hce5: data = 9'o0;
		14'hce6: data = 9'o0;
		14'hce7: data = 9'o0;
		14'hce8: data = 9'o0;
		14'hce9: data = 9'o0;
		14'hcea: data = 9'o0;
		14'hceb: data = 9'o541;
		14'hcec: data = 9'o762;
		14'hced: data = 9'o773;
		14'hcee: data = 9'o252;
		14'hcef: data = 9'o52;
		14'hcf0: data = 9'o52;
		14'hcf1: data = 9'o52;
		14'hcf2: data = 9'o152;
		14'hcf3: data = 9'o142;
		14'hcf4: data = 9'o242;
		14'hcf5: data = 9'o142;
		14'hcf6: data = 9'o152;
		14'hcf7: data = 9'o152;
		14'hcf8: data = 9'o152;
		14'hcf9: data = 9'o142;
		14'hcfa: data = 9'o142;
		14'hcfb: data = 9'o152;
		14'hcfc: data = 9'o52;
		14'hcfd: data = 9'o52;
		14'hcfe: data = 9'o152;
		14'hcff: data = 9'o142;
		14'hd00: data = 9'o142;
		14'hd01: data = 9'o142;
		14'hd02: data = 9'o153;
		14'hd03: data = 9'o52;
		14'hd04: data = 9'o52;
		14'hd05: data = 9'o152;
		14'hd06: data = 9'o573;
		14'hd07: data = 9'o773;
		14'hd08: data = 9'o773;
		14'hd09: data = 9'o773;
		14'hd0a: data = 9'o773;
		14'hd0b: data = 9'o773;
		14'hd0c: data = 9'o773;
		14'hd0d: data = 9'o773;
		14'hd0e: data = 9'o773;
		14'hd0f: data = 9'o773;
		14'hd10: data = 9'o773;
		14'hd11: data = 9'o463;
		14'hd12: data = 9'o152;
		14'hd13: data = 9'o152;
		14'hd14: data = 9'o52;
		14'hd15: data = 9'o152;
		14'hd16: data = 9'o152;
		14'hd17: data = 9'o152;
		14'hd18: data = 9'o363;
		14'hd19: data = 9'o773;
		14'hd1a: data = 9'o773;
		14'hd1b: data = 9'o773;
		14'hd1c: data = 9'o773;
		14'hd1d: data = 9'o773;
		14'hd1e: data = 9'o773;
		14'hd1f: data = 9'o773;
		14'hd20: data = 9'o773;
		14'hd21: data = 9'o773;
		14'hd22: data = 9'o773;
		14'hd23: data = 9'o673;
		14'hd24: data = 9'o152;
		14'hd25: data = 9'o152;
		14'hd26: data = 9'o52;
		14'hd27: data = 9'o152;
		14'hd28: data = 9'o152;
		14'hd29: data = 9'o252;
		14'hd2a: data = 9'o142;
		14'hd2b: data = 9'o142;
		14'hd2c: data = 9'o152;
		14'hd2d: data = 9'o152;
		14'hd2e: data = 9'o152;
		14'hd2f: data = 9'o152;
		14'hd30: data = 9'o152;
		14'hd31: data = 9'o152;
		14'hd32: data = 9'o152;
		14'hd33: data = 9'o152;
		14'hd34: data = 9'o152;
		14'hd35: data = 9'o142;
		14'hd36: data = 9'o242;
		14'hd37: data = 9'o142;
		14'hd38: data = 9'o152;
		14'hd39: data = 9'o52;
		14'hd3a: data = 9'o152;
		14'hd3b: data = 9'o252;
		14'hd3c: data = 9'o773;
		14'hd3d: data = 9'o662;
		14'hd3e: data = 9'o0;
		14'hd3f: data = 9'o0;
		14'hd40: data = 9'o0;
		14'hd41: data = 9'o0;
		14'hd42: data = 9'o0;
		14'hd43: data = 9'o0;
		14'hd44: data = 9'o0;
		14'hd45: data = 9'o0;
		14'hd46: data = 9'o0;
		14'hd47: data = 9'o0;
		14'hd48: data = 9'o0;
		14'hd49: data = 9'o0;
		14'hd4a: data = 9'o0;
		14'hd4b: data = 9'o0;
		14'hd4c: data = 9'o0;
		14'hd4d: data = 9'o0;
		14'hd4e: data = 9'o0;
		14'hd4f: data = 9'o551;
		14'hd50: data = 9'o662;
		14'hd51: data = 9'o673;
		14'hd52: data = 9'o252;
		14'hd53: data = 9'o152;
		14'hd54: data = 9'o52;
		14'hd55: data = 9'o52;
		14'hd56: data = 9'o52;
		14'hd57: data = 9'o152;
		14'hd58: data = 9'o152;
		14'hd59: data = 9'o152;
		14'hd5a: data = 9'o152;
		14'hd5b: data = 9'o52;
		14'hd5c: data = 9'o152;
		14'hd5d: data = 9'o152;
		14'hd5e: data = 9'o152;
		14'hd5f: data = 9'o152;
		14'hd60: data = 9'o52;
		14'hd61: data = 9'o53;
		14'hd62: data = 9'o52;
		14'hd63: data = 9'o152;
		14'hd64: data = 9'o152;
		14'hd65: data = 9'o152;
		14'hd66: data = 9'o152;
		14'hd67: data = 9'o152;
		14'hd68: data = 9'o152;
		14'hd69: data = 9'o152;
		14'hd6a: data = 9'o573;
		14'hd6b: data = 9'o773;
		14'hd6c: data = 9'o773;
		14'hd6d: data = 9'o773;
		14'hd6e: data = 9'o773;
		14'hd6f: data = 9'o773;
		14'hd70: data = 9'o773;
		14'hd71: data = 9'o773;
		14'hd72: data = 9'o773;
		14'hd73: data = 9'o773;
		14'hd74: data = 9'o773;
		14'hd75: data = 9'o352;
		14'hd76: data = 9'o152;
		14'hd77: data = 9'o152;
		14'hd78: data = 9'o152;
		14'hd79: data = 9'o152;
		14'hd7a: data = 9'o52;
		14'hd7b: data = 9'o152;
		14'hd7c: data = 9'o352;
		14'hd7d: data = 9'o673;
		14'hd7e: data = 9'o773;
		14'hd7f: data = 9'o773;
		14'hd80: data = 9'o773;
		14'hd81: data = 9'o773;
		14'hd82: data = 9'o773;
		14'hd83: data = 9'o773;
		14'hd84: data = 9'o773;
		14'hd85: data = 9'o773;
		14'hd86: data = 9'o773;
		14'hd87: data = 9'o573;
		14'hd88: data = 9'o152;
		14'hd89: data = 9'o152;
		14'hd8a: data = 9'o152;
		14'hd8b: data = 9'o52;
		14'hd8c: data = 9'o152;
		14'hd8d: data = 9'o152;
		14'hd8e: data = 9'o152;
		14'hd8f: data = 9'o152;
		14'hd90: data = 9'o152;
		14'hd91: data = 9'o152;
		14'hd92: data = 9'o152;
		14'hd93: data = 9'o152;
		14'hd94: data = 9'o152;
		14'hd95: data = 9'o152;
		14'hd96: data = 9'o152;
		14'hd97: data = 9'o152;
		14'hd98: data = 9'o152;
		14'hd99: data = 9'o152;
		14'hd9a: data = 9'o152;
		14'hd9b: data = 9'o152;
		14'hd9c: data = 9'o52;
		14'hd9d: data = 9'o152;
		14'hd9e: data = 9'o152;
		14'hd9f: data = 9'o252;
		14'hda0: data = 9'o773;
		14'hda1: data = 9'o763;
		14'hda2: data = 9'o0;
		14'hda3: data = 9'o0;
		14'hda4: data = 9'o0;
		14'hda5: data = 9'o0;
		14'hda6: data = 9'o0;
		14'hda7: data = 9'o0;
		14'hda8: data = 9'o0;
		14'hda9: data = 9'o0;
		14'hdaa: data = 9'o0;
		14'hdab: data = 9'o0;
		14'hdac: data = 9'o0;
		14'hdad: data = 9'o0;
		14'hdae: data = 9'o0;
		14'hdaf: data = 9'o0;
		14'hdb0: data = 9'o0;
		14'hdb1: data = 9'o0;
		14'hdb2: data = 9'o0;
		14'hdb3: data = 9'o551;
		14'hdb4: data = 9'o663;
		14'hdb5: data = 9'o773;
		14'hdb6: data = 9'o252;
		14'hdb7: data = 9'o152;
		14'hdb8: data = 9'o152;
		14'hdb9: data = 9'o52;
		14'hdba: data = 9'o52;
		14'hdbb: data = 9'o52;
		14'hdbc: data = 9'o152;
		14'hdbd: data = 9'o152;
		14'hdbe: data = 9'o52;
		14'hdbf: data = 9'o52;
		14'hdc0: data = 9'o52;
		14'hdc1: data = 9'o52;
		14'hdc2: data = 9'o52;
		14'hdc3: data = 9'o52;
		14'hdc4: data = 9'o52;
		14'hdc5: data = 9'o52;
		14'hdc6: data = 9'o52;
		14'hdc7: data = 9'o52;
		14'hdc8: data = 9'o52;
		14'hdc9: data = 9'o152;
		14'hdca: data = 9'o152;
		14'hdcb: data = 9'o142;
		14'hdcc: data = 9'o152;
		14'hdcd: data = 9'o152;
		14'hdce: data = 9'o573;
		14'hdcf: data = 9'o773;
		14'hdd0: data = 9'o773;
		14'hdd1: data = 9'o773;
		14'hdd2: data = 9'o773;
		14'hdd3: data = 9'o773;
		14'hdd4: data = 9'o773;
		14'hdd5: data = 9'o773;
		14'hdd6: data = 9'o773;
		14'hdd7: data = 9'o773;
		14'hdd8: data = 9'o673;
		14'hdd9: data = 9'o252;
		14'hdda: data = 9'o152;
		14'hddb: data = 9'o152;
		14'hddc: data = 9'o152;
		14'hddd: data = 9'o152;
		14'hdde: data = 9'o52;
		14'hddf: data = 9'o152;
		14'hde0: data = 9'o252;
		14'hde1: data = 9'o673;
		14'hde2: data = 9'o773;
		14'hde3: data = 9'o773;
		14'hde4: data = 9'o773;
		14'hde5: data = 9'o773;
		14'hde6: data = 9'o773;
		14'hde7: data = 9'o773;
		14'hde8: data = 9'o773;
		14'hde9: data = 9'o773;
		14'hdea: data = 9'o773;
		14'hdeb: data = 9'o673;
		14'hdec: data = 9'o142;
		14'hded: data = 9'o152;
		14'hdee: data = 9'o52;
		14'hdef: data = 9'o52;
		14'hdf0: data = 9'o152;
		14'hdf1: data = 9'o152;
		14'hdf2: data = 9'o152;
		14'hdf3: data = 9'o152;
		14'hdf4: data = 9'o152;
		14'hdf5: data = 9'o52;
		14'hdf6: data = 9'o152;
		14'hdf7: data = 9'o152;
		14'hdf8: data = 9'o152;
		14'hdf9: data = 9'o52;
		14'hdfa: data = 9'o52;
		14'hdfb: data = 9'o52;
		14'hdfc: data = 9'o52;
		14'hdfd: data = 9'o52;
		14'hdfe: data = 9'o152;
		14'hdff: data = 9'o152;
		14'he00: data = 9'o152;
		14'he01: data = 9'o152;
		14'he02: data = 9'o152;
		14'he03: data = 9'o252;
		14'he04: data = 9'o773;
		14'he05: data = 9'o662;
		14'he06: data = 9'o0;
		14'he07: data = 9'o0;
		14'he08: data = 9'o0;
		14'he09: data = 9'o0;
		14'he0a: data = 9'o0;
		14'he0b: data = 9'o0;
		14'he0c: data = 9'o0;
		14'he0d: data = 9'o0;
		14'he0e: data = 9'o0;
		14'he0f: data = 9'o0;
		14'he10: data = 9'o0;
		14'he11: data = 9'o0;
		14'he12: data = 9'o0;
		14'he13: data = 9'o0;
		14'he14: data = 9'o0;
		14'he15: data = 9'o0;
		14'he16: data = 9'o0;
		14'he17: data = 9'o551;
		14'he18: data = 9'o663;
		14'he19: data = 9'o773;
		14'he1a: data = 9'o352;
		14'he1b: data = 9'o142;
		14'he1c: data = 9'o152;
		14'he1d: data = 9'o152;
		14'he1e: data = 9'o52;
		14'he1f: data = 9'o52;
		14'he20: data = 9'o52;
		14'he21: data = 9'o152;
		14'he22: data = 9'o52;
		14'he23: data = 9'o52;
		14'he24: data = 9'o52;
		14'he25: data = 9'o52;
		14'he26: data = 9'o52;
		14'he27: data = 9'o52;
		14'he28: data = 9'o52;
		14'he29: data = 9'o52;
		14'he2a: data = 9'o52;
		14'he2b: data = 9'o52;
		14'he2c: data = 9'o52;
		14'he2d: data = 9'o152;
		14'he2e: data = 9'o252;
		14'he2f: data = 9'o142;
		14'he30: data = 9'o152;
		14'he31: data = 9'o252;
		14'he32: data = 9'o573;
		14'he33: data = 9'o773;
		14'he34: data = 9'o773;
		14'he35: data = 9'o773;
		14'he36: data = 9'o773;
		14'he37: data = 9'o673;
		14'he38: data = 9'o673;
		14'he39: data = 9'o673;
		14'he3a: data = 9'o773;
		14'he3b: data = 9'o773;
		14'he3c: data = 9'o573;
		14'he3d: data = 9'o252;
		14'he3e: data = 9'o152;
		14'he3f: data = 9'o152;
		14'he40: data = 9'o152;
		14'he41: data = 9'o52;
		14'he42: data = 9'o52;
		14'he43: data = 9'o152;
		14'he44: data = 9'o152;
		14'he45: data = 9'o573;
		14'he46: data = 9'o773;
		14'he47: data = 9'o773;
		14'he48: data = 9'o673;
		14'he49: data = 9'o673;
		14'he4a: data = 9'o673;
		14'he4b: data = 9'o773;
		14'he4c: data = 9'o773;
		14'he4d: data = 9'o773;
		14'he4e: data = 9'o773;
		14'he4f: data = 9'o673;
		14'he50: data = 9'o242;
		14'he51: data = 9'o152;
		14'he52: data = 9'o152;
		14'he53: data = 9'o152;
		14'he54: data = 9'o152;
		14'he55: data = 9'o52;
		14'he56: data = 9'o52;
		14'he57: data = 9'o52;
		14'he58: data = 9'o52;
		14'he59: data = 9'o52;
		14'he5a: data = 9'o52;
		14'he5b: data = 9'o52;
		14'he5c: data = 9'o52;
		14'he5d: data = 9'o52;
		14'he5e: data = 9'o52;
		14'he5f: data = 9'o52;
		14'he60: data = 9'o52;
		14'he61: data = 9'o52;
		14'he62: data = 9'o52;
		14'he63: data = 9'o152;
		14'he64: data = 9'o152;
		14'he65: data = 9'o142;
		14'he66: data = 9'o152;
		14'he67: data = 9'o352;
		14'he68: data = 9'o773;
		14'he69: data = 9'o762;
		14'he6a: data = 9'o0;
		14'he6b: data = 9'o0;
		14'he6c: data = 9'o0;
		14'he6d: data = 9'o0;
		14'he6e: data = 9'o0;
		14'he6f: data = 9'o0;
		14'he70: data = 9'o0;
		14'he71: data = 9'o0;
		14'he72: data = 9'o0;
		14'he73: data = 9'o0;
		14'he74: data = 9'o0;
		14'he75: data = 9'o0;
		14'he76: data = 9'o0;
		14'he77: data = 9'o0;
		14'he78: data = 9'o0;
		14'he79: data = 9'o0;
		14'he7a: data = 9'o0;
		14'he7b: data = 9'o652;
		14'he7c: data = 9'o662;
		14'he7d: data = 9'o773;
		14'he7e: data = 9'o352;
		14'he7f: data = 9'o242;
		14'he80: data = 9'o242;
		14'he81: data = 9'o152;
		14'he82: data = 9'o152;
		14'he83: data = 9'o52;
		14'he84: data = 9'o52;
		14'he85: data = 9'o52;
		14'he86: data = 9'o52;
		14'he87: data = 9'o52;
		14'he88: data = 9'o52;
		14'he89: data = 9'o52;
		14'he8a: data = 9'o52;
		14'he8b: data = 9'o52;
		14'he8c: data = 9'o52;
		14'he8d: data = 9'o52;
		14'he8e: data = 9'o52;
		14'he8f: data = 9'o152;
		14'he90: data = 9'o52;
		14'he91: data = 9'o152;
		14'he92: data = 9'o242;
		14'he93: data = 9'o242;
		14'he94: data = 9'o242;
		14'he95: data = 9'o352;
		14'he96: data = 9'o673;
		14'he97: data = 9'o773;
		14'he98: data = 9'o773;
		14'he99: data = 9'o773;
		14'he9a: data = 9'o463;
		14'he9b: data = 9'o242;
		14'he9c: data = 9'o252;
		14'he9d: data = 9'o352;
		14'he9e: data = 9'o673;
		14'he9f: data = 9'o773;
		14'hea0: data = 9'o463;
		14'hea1: data = 9'o152;
		14'hea2: data = 9'o152;
		14'hea3: data = 9'o152;
		14'hea4: data = 9'o152;
		14'hea5: data = 9'o52;
		14'hea6: data = 9'o52;
		14'hea7: data = 9'o152;
		14'hea8: data = 9'o142;
		14'hea9: data = 9'o463;
		14'heaa: data = 9'o773;
		14'heab: data = 9'o673;
		14'heac: data = 9'o252;
		14'head: data = 9'o152;
		14'heae: data = 9'o252;
		14'heaf: data = 9'o463;
		14'heb0: data = 9'o673;
		14'heb1: data = 9'o773;
		14'heb2: data = 9'o773;
		14'heb3: data = 9'o673;
		14'heb4: data = 9'o342;
		14'heb5: data = 9'o242;
		14'heb6: data = 9'o142;
		14'heb7: data = 9'o152;
		14'heb8: data = 9'o52;
		14'heb9: data = 9'o52;
		14'heba: data = 9'o52;
		14'hebb: data = 9'o52;
		14'hebc: data = 9'o52;
		14'hebd: data = 9'o52;
		14'hebe: data = 9'o52;
		14'hebf: data = 9'o52;
		14'hec0: data = 9'o52;
		14'hec1: data = 9'o52;
		14'hec2: data = 9'o52;
		14'hec3: data = 9'o52;
		14'hec4: data = 9'o52;
		14'hec5: data = 9'o52;
		14'hec6: data = 9'o52;
		14'hec7: data = 9'o152;
		14'hec8: data = 9'o252;
		14'hec9: data = 9'o242;
		14'heca: data = 9'o242;
		14'hecb: data = 9'o352;
		14'hecc: data = 9'o773;
		14'hecd: data = 9'o762;
		14'hece: data = 9'o0;
		14'hecf: data = 9'o0;
		14'hed0: data = 9'o0;
		14'hed1: data = 9'o0;
		14'hed2: data = 9'o0;
		14'hed3: data = 9'o0;
		14'hed4: data = 9'o0;
		14'hed5: data = 9'o0;
		14'hed6: data = 9'o0;
		14'hed7: data = 9'o0;
		14'hed8: data = 9'o0;
		14'hed9: data = 9'o0;
		14'heda: data = 9'o0;
		14'hedb: data = 9'o0;
		14'hedc: data = 9'o0;
		14'hedd: data = 9'o0;
		14'hede: data = 9'o0;
		14'hedf: data = 9'o651;
		14'hee0: data = 9'o662;
		14'hee1: data = 9'o773;
		14'hee2: data = 9'o673;
		14'hee3: data = 9'o673;
		14'hee4: data = 9'o673;
		14'hee5: data = 9'o573;
		14'hee6: data = 9'o373;
		14'hee7: data = 9'o273;
		14'hee8: data = 9'o172;
		14'hee9: data = 9'o172;
		14'heea: data = 9'o172;
		14'heeb: data = 9'o173;
		14'heec: data = 9'o273;
		14'heed: data = 9'o272;
		14'heee: data = 9'o272;
		14'heef: data = 9'o172;
		14'hef0: data = 9'o173;
		14'hef1: data = 9'o173;
		14'hef2: data = 9'o272;
		14'hef3: data = 9'o272;
		14'hef4: data = 9'o272;
		14'hef5: data = 9'o272;
		14'hef6: data = 9'o573;
		14'hef7: data = 9'o673;
		14'hef8: data = 9'o573;
		14'hef9: data = 9'o673;
		14'hefa: data = 9'o773;
		14'hefb: data = 9'o773;
		14'hefc: data = 9'o773;
		14'hefd: data = 9'o773;
		14'hefe: data = 9'o463;
		14'heff: data = 9'o142;
		14'hf00: data = 9'o152;
		14'hf01: data = 9'o242;
		14'hf02: data = 9'o673;
		14'hf03: data = 9'o773;
		14'hf04: data = 9'o362;
		14'hf05: data = 9'o152;
		14'hf06: data = 9'o152;
		14'hf07: data = 9'o152;
		14'hf08: data = 9'o52;
		14'hf09: data = 9'o52;
		14'hf0a: data = 9'o52;
		14'hf0b: data = 9'o152;
		14'hf0c: data = 9'o142;
		14'hf0d: data = 9'o363;
		14'hf0e: data = 9'o673;
		14'hf0f: data = 9'o673;
		14'hf10: data = 9'o152;
		14'hf11: data = 9'o152;
		14'hf12: data = 9'o152;
		14'hf13: data = 9'o363;
		14'hf14: data = 9'o673;
		14'hf15: data = 9'o773;
		14'hf16: data = 9'o773;
		14'hf17: data = 9'o773;
		14'hf18: data = 9'o673;
		14'hf19: data = 9'o673;
		14'hf1a: data = 9'o673;
		14'hf1b: data = 9'o573;
		14'hf1c: data = 9'o273;
		14'hf1d: data = 9'o173;
		14'hf1e: data = 9'o172;
		14'hf1f: data = 9'o172;
		14'hf20: data = 9'o173;
		14'hf21: data = 9'o173;
		14'hf22: data = 9'o173;
		14'hf23: data = 9'o172;
		14'hf24: data = 9'o172;
		14'hf25: data = 9'o272;
		14'hf26: data = 9'o273;
		14'hf27: data = 9'o273;
		14'hf28: data = 9'o173;
		14'hf29: data = 9'o172;
		14'hf2a: data = 9'o272;
		14'hf2b: data = 9'o373;
		14'hf2c: data = 9'o573;
		14'hf2d: data = 9'o673;
		14'hf2e: data = 9'o673;
		14'hf2f: data = 9'o673;
		14'hf30: data = 9'o773;
		14'hf31: data = 9'o773;
		14'hf32: data = 9'o0;
		14'hf33: data = 9'o0;
		14'hf34: data = 9'o0;
		14'hf35: data = 9'o0;
		14'hf36: data = 9'o0;
		14'hf37: data = 9'o0;
		14'hf38: data = 9'o0;
		14'hf39: data = 9'o0;
		14'hf3a: data = 9'o0;
		14'hf3b: data = 9'o0;
		14'hf3c: data = 9'o0;
		14'hf3d: data = 9'o0;
		14'hf3e: data = 9'o0;
		14'hf3f: data = 9'o0;
		14'hf40: data = 9'o0;
		14'hf41: data = 9'o0;
		14'hf42: data = 9'o0;
		14'hf43: data = 9'o651;
		14'hf44: data = 9'o662;
		14'hf45: data = 9'o773;
		14'hf46: data = 9'o773;
		14'hf47: data = 9'o773;
		14'hf48: data = 9'o773;
		14'hf49: data = 9'o673;
		14'hf4a: data = 9'o473;
		14'hf4b: data = 9'o273;
		14'hf4c: data = 9'o272;
		14'hf4d: data = 9'o172;
		14'hf4e: data = 9'o172;
		14'hf4f: data = 9'o272;
		14'hf50: data = 9'o273;
		14'hf51: data = 9'o272;
		14'hf52: data = 9'o272;
		14'hf53: data = 9'o272;
		14'hf54: data = 9'o272;
		14'hf55: data = 9'o273;
		14'hf56: data = 9'o272;
		14'hf57: data = 9'o272;
		14'hf58: data = 9'o172;
		14'hf59: data = 9'o272;
		14'hf5a: data = 9'o573;
		14'hf5b: data = 9'o773;
		14'hf5c: data = 9'o773;
		14'hf5d: data = 9'o773;
		14'hf5e: data = 9'o773;
		14'hf5f: data = 9'o773;
		14'hf60: data = 9'o773;
		14'hf61: data = 9'o773;
		14'hf62: data = 9'o463;
		14'hf63: data = 9'o152;
		14'hf64: data = 9'o152;
		14'hf65: data = 9'o252;
		14'hf66: data = 9'o673;
		14'hf67: data = 9'o673;
		14'hf68: data = 9'o252;
		14'hf69: data = 9'o152;
		14'hf6a: data = 9'o152;
		14'hf6b: data = 9'o152;
		14'hf6c: data = 9'o52;
		14'hf6d: data = 9'o52;
		14'hf6e: data = 9'o52;
		14'hf6f: data = 9'o152;
		14'hf70: data = 9'o152;
		14'hf71: data = 9'o252;
		14'hf72: data = 9'o673;
		14'hf73: data = 9'o673;
		14'hf74: data = 9'o252;
		14'hf75: data = 9'o152;
		14'hf76: data = 9'o242;
		14'hf77: data = 9'o463;
		14'hf78: data = 9'o773;
		14'hf79: data = 9'o773;
		14'hf7a: data = 9'o773;
		14'hf7b: data = 9'o773;
		14'hf7c: data = 9'o773;
		14'hf7d: data = 9'o773;
		14'hf7e: data = 9'o773;
		14'hf7f: data = 9'o673;
		14'hf80: data = 9'o373;
		14'hf81: data = 9'o273;
		14'hf82: data = 9'o172;
		14'hf83: data = 9'o172;
		14'hf84: data = 9'o173;
		14'hf85: data = 9'o173;
		14'hf86: data = 9'o173;
		14'hf87: data = 9'o172;
		14'hf88: data = 9'o272;
		14'hf89: data = 9'o272;
		14'hf8a: data = 9'o273;
		14'hf8b: data = 9'o273;
		14'hf8c: data = 9'o273;
		14'hf8d: data = 9'o272;
		14'hf8e: data = 9'o272;
		14'hf8f: data = 9'o473;
		14'hf90: data = 9'o673;
		14'hf91: data = 9'o773;
		14'hf92: data = 9'o773;
		14'hf93: data = 9'o773;
		14'hf94: data = 9'o773;
		14'hf95: data = 9'o762;
		14'hf96: data = 9'o0;
		14'hf97: data = 9'o0;
		14'hf98: data = 9'o0;
		14'hf99: data = 9'o0;
		14'hf9a: data = 9'o0;
		14'hf9b: data = 9'o0;
		14'hf9c: data = 9'o0;
		14'hf9d: data = 9'o0;
		14'hf9e: data = 9'o0;
		14'hf9f: data = 9'o0;
		14'hfa0: data = 9'o0;
		14'hfa1: data = 9'o0;
		14'hfa2: data = 9'o0;
		14'hfa3: data = 9'o0;
		14'hfa4: data = 9'o0;
		14'hfa5: data = 9'o0;
		14'hfa6: data = 9'o0;
		14'hfa7: data = 9'o652;
		14'hfa8: data = 9'o662;
		14'hfa9: data = 9'o773;
		14'hfaa: data = 9'o773;
		14'hfab: data = 9'o773;
		14'hfac: data = 9'o773;
		14'hfad: data = 9'o773;
		14'hfae: data = 9'o373;
		14'hfaf: data = 9'o272;
		14'hfb0: data = 9'o172;
		14'hfb1: data = 9'o172;
		14'hfb2: data = 9'o172;
		14'hfb3: data = 9'o172;
		14'hfb4: data = 9'o272;
		14'hfb5: data = 9'o272;
		14'hfb6: data = 9'o272;
		14'hfb7: data = 9'o272;
		14'hfb8: data = 9'o172;
		14'hfb9: data = 9'o172;
		14'hfba: data = 9'o272;
		14'hfbb: data = 9'o272;
		14'hfbc: data = 9'o172;
		14'hfbd: data = 9'o272;
		14'hfbe: data = 9'o573;
		14'hfbf: data = 9'o773;
		14'hfc0: data = 9'o773;
		14'hfc1: data = 9'o773;
		14'hfc2: data = 9'o773;
		14'hfc3: data = 9'o773;
		14'hfc4: data = 9'o773;
		14'hfc5: data = 9'o773;
		14'hfc6: data = 9'o463;
		14'hfc7: data = 9'o152;
		14'hfc8: data = 9'o152;
		14'hfc9: data = 9'o152;
		14'hfca: data = 9'o573;
		14'hfcb: data = 9'o573;
		14'hfcc: data = 9'o152;
		14'hfcd: data = 9'o52;
		14'hfce: data = 9'o152;
		14'hfcf: data = 9'o152;
		14'hfd0: data = 9'o52;
		14'hfd1: data = 9'o52;
		14'hfd2: data = 9'o52;
		14'hfd3: data = 9'o152;
		14'hfd4: data = 9'o152;
		14'hfd5: data = 9'o252;
		14'hfd6: data = 9'o573;
		14'hfd7: data = 9'o573;
		14'hfd8: data = 9'o152;
		14'hfd9: data = 9'o152;
		14'hfda: data = 9'o142;
		14'hfdb: data = 9'o463;
		14'hfdc: data = 9'o773;
		14'hfdd: data = 9'o773;
		14'hfde: data = 9'o773;
		14'hfdf: data = 9'o773;
		14'hfe0: data = 9'o773;
		14'hfe1: data = 9'o773;
		14'hfe2: data = 9'o773;
		14'hfe3: data = 9'o673;
		14'hfe4: data = 9'o272;
		14'hfe5: data = 9'o272;
		14'hfe6: data = 9'o172;
		14'hfe7: data = 9'o172;
		14'hfe8: data = 9'o172;
		14'hfe9: data = 9'o173;
		14'hfea: data = 9'o172;
		14'hfeb: data = 9'o172;
		14'hfec: data = 9'o272;
		14'hfed: data = 9'o272;
		14'hfee: data = 9'o273;
		14'hfef: data = 9'o272;
		14'hff0: data = 9'o273;
		14'hff1: data = 9'o172;
		14'hff2: data = 9'o272;
		14'hff3: data = 9'o373;
		14'hff4: data = 9'o673;
		14'hff5: data = 9'o773;
		14'hff6: data = 9'o773;
		14'hff7: data = 9'o773;
		14'hff8: data = 9'o773;
		14'hff9: data = 9'o662;
		14'hffa: data = 9'o0;
		14'hffb: data = 9'o0;
		14'hffc: data = 9'o0;
		14'hffd: data = 9'o0;
		14'hffe: data = 9'o0;
		14'hfff: data = 9'o0;
		14'h1000: data = 9'o0;
		14'h1001: data = 9'o0;
		14'h1002: data = 9'o0;
		14'h1003: data = 9'o0;
		14'h1004: data = 9'o0;
		14'h1005: data = 9'o0;
		14'h1006: data = 9'o0;
		14'h1007: data = 9'o0;
		14'h1008: data = 9'o0;
		14'h1009: data = 9'o0;
		14'h100a: data = 9'o0;
		14'h100b: data = 9'o652;
		14'h100c: data = 9'o662;
		14'h100d: data = 9'o773;
		14'h100e: data = 9'o773;
		14'h100f: data = 9'o773;
		14'h1010: data = 9'o773;
		14'h1011: data = 9'o673;
		14'h1012: data = 9'o372;
		14'h1013: data = 9'o272;
		14'h1014: data = 9'o172;
		14'h1015: data = 9'o172;
		14'h1016: data = 9'o172;
		14'h1017: data = 9'o173;
		14'h1018: data = 9'o172;
		14'h1019: data = 9'o172;
		14'h101a: data = 9'o272;
		14'h101b: data = 9'o172;
		14'h101c: data = 9'o172;
		14'h101d: data = 9'o172;
		14'h101e: data = 9'o272;
		14'h101f: data = 9'o272;
		14'h1020: data = 9'o172;
		14'h1021: data = 9'o272;
		14'h1022: data = 9'o573;
		14'h1023: data = 9'o773;
		14'h1024: data = 9'o773;
		14'h1025: data = 9'o773;
		14'h1026: data = 9'o773;
		14'h1027: data = 9'o773;
		14'h1028: data = 9'o773;
		14'h1029: data = 9'o773;
		14'h102a: data = 9'o463;
		14'h102b: data = 9'o152;
		14'h102c: data = 9'o152;
		14'h102d: data = 9'o152;
		14'h102e: data = 9'o253;
		14'h102f: data = 9'o252;
		14'h1030: data = 9'o152;
		14'h1031: data = 9'o52;
		14'h1032: data = 9'o52;
		14'h1033: data = 9'o52;
		14'h1034: data = 9'o52;
		14'h1035: data = 9'o52;
		14'h1036: data = 9'o52;
		14'h1037: data = 9'o52;
		14'h1038: data = 9'o152;
		14'h1039: data = 9'o152;
		14'h103a: data = 9'o152;
		14'h103b: data = 9'o152;
		14'h103c: data = 9'o152;
		14'h103d: data = 9'o152;
		14'h103e: data = 9'o152;
		14'h103f: data = 9'o363;
		14'h1040: data = 9'o773;
		14'h1041: data = 9'o773;
		14'h1042: data = 9'o773;
		14'h1043: data = 9'o773;
		14'h1044: data = 9'o773;
		14'h1045: data = 9'o773;
		14'h1046: data = 9'o673;
		14'h1047: data = 9'o573;
		14'h1048: data = 9'o272;
		14'h1049: data = 9'o272;
		14'h104a: data = 9'o172;
		14'h104b: data = 9'o172;
		14'h104c: data = 9'o172;
		14'h104d: data = 9'o172;
		14'h104e: data = 9'o172;
		14'h104f: data = 9'o272;
		14'h1050: data = 9'o272;
		14'h1051: data = 9'o272;
		14'h1052: data = 9'o272;
		14'h1053: data = 9'o273;
		14'h1054: data = 9'o172;
		14'h1055: data = 9'o172;
		14'h1056: data = 9'o272;
		14'h1057: data = 9'o372;
		14'h1058: data = 9'o673;
		14'h1059: data = 9'o773;
		14'h105a: data = 9'o773;
		14'h105b: data = 9'o773;
		14'h105c: data = 9'o773;
		14'h105d: data = 9'o662;
		14'h105e: data = 9'o0;
		14'h105f: data = 9'o0;
		14'h1060: data = 9'o0;
		14'h1061: data = 9'o0;
		14'h1062: data = 9'o0;
		14'h1063: data = 9'o0;
		14'h1064: data = 9'o0;
		14'h1065: data = 9'o0;
		14'h1066: data = 9'o0;
		14'h1067: data = 9'o0;
		14'h1068: data = 9'o0;
		14'h1069: data = 9'o0;
		14'h106a: data = 9'o0;
		14'h106b: data = 9'o0;
		14'h106c: data = 9'o0;
		14'h106d: data = 9'o0;
		14'h106e: data = 9'o0;
		14'h106f: data = 9'o652;
		14'h1070: data = 9'o662;
		14'h1071: data = 9'o773;
		14'h1072: data = 9'o773;
		14'h1073: data = 9'o773;
		14'h1074: data = 9'o773;
		14'h1075: data = 9'o673;
		14'h1076: data = 9'o372;
		14'h1077: data = 9'o272;
		14'h1078: data = 9'o172;
		14'h1079: data = 9'o172;
		14'h107a: data = 9'o172;
		14'h107b: data = 9'o172;
		14'h107c: data = 9'o273;
		14'h107d: data = 9'o272;
		14'h107e: data = 9'o272;
		14'h107f: data = 9'o272;
		14'h1080: data = 9'o273;
		14'h1081: data = 9'o172;
		14'h1082: data = 9'o172;
		14'h1083: data = 9'o172;
		14'h1084: data = 9'o172;
		14'h1085: data = 9'o272;
		14'h1086: data = 9'o473;
		14'h1087: data = 9'o773;
		14'h1088: data = 9'o773;
		14'h1089: data = 9'o773;
		14'h108a: data = 9'o773;
		14'h108b: data = 9'o773;
		14'h108c: data = 9'o773;
		14'h108d: data = 9'o773;
		14'h108e: data = 9'o463;
		14'h108f: data = 9'o152;
		14'h1090: data = 9'o152;
		14'h1091: data = 9'o152;
		14'h1092: data = 9'o152;
		14'h1093: data = 9'o152;
		14'h1094: data = 9'o152;
		14'h1095: data = 9'o52;
		14'h1096: data = 9'o52;
		14'h1097: data = 9'o52;
		14'h1098: data = 9'o152;
		14'h1099: data = 9'o152;
		14'h109a: data = 9'o52;
		14'h109b: data = 9'o52;
		14'h109c: data = 9'o152;
		14'h109d: data = 9'o152;
		14'h109e: data = 9'o52;
		14'h109f: data = 9'o52;
		14'h10a0: data = 9'o152;
		14'h10a1: data = 9'o152;
		14'h10a2: data = 9'o152;
		14'h10a3: data = 9'o363;
		14'h10a4: data = 9'o773;
		14'h10a5: data = 9'o773;
		14'h10a6: data = 9'o773;
		14'h10a7: data = 9'o773;
		14'h10a8: data = 9'o773;
		14'h10a9: data = 9'o773;
		14'h10aa: data = 9'o673;
		14'h10ab: data = 9'o473;
		14'h10ac: data = 9'o272;
		14'h10ad: data = 9'o272;
		14'h10ae: data = 9'o272;
		14'h10af: data = 9'o172;
		14'h10b0: data = 9'o172;
		14'h10b1: data = 9'o272;
		14'h10b2: data = 9'o272;
		14'h10b3: data = 9'o272;
		14'h10b4: data = 9'o272;
		14'h10b5: data = 9'o272;
		14'h10b6: data = 9'o272;
		14'h10b7: data = 9'o172;
		14'h10b8: data = 9'o172;
		14'h10b9: data = 9'o172;
		14'h10ba: data = 9'o172;
		14'h10bb: data = 9'o372;
		14'h10bc: data = 9'o673;
		14'h10bd: data = 9'o773;
		14'h10be: data = 9'o773;
		14'h10bf: data = 9'o773;
		14'h10c0: data = 9'o773;
		14'h10c1: data = 9'o662;
		14'h10c2: data = 9'o0;
		14'h10c3: data = 9'o0;
		14'h10c4: data = 9'o0;
		14'h10c5: data = 9'o0;
		14'h10c6: data = 9'o0;
		14'h10c7: data = 9'o0;
		14'h10c8: data = 9'o0;
		14'h10c9: data = 9'o0;
		14'h10ca: data = 9'o0;
		14'h10cb: data = 9'o0;
		14'h10cc: data = 9'o0;
		14'h10cd: data = 9'o0;
		14'h10ce: data = 9'o0;
		14'h10cf: data = 9'o0;
		14'h10d0: data = 9'o0;
		14'h10d1: data = 9'o0;
		14'h10d2: data = 9'o0;
		14'h10d3: data = 9'o652;
		14'h10d4: data = 9'o762;
		14'h10d5: data = 9'o773;
		14'h10d6: data = 9'o773;
		14'h10d7: data = 9'o773;
		14'h10d8: data = 9'o773;
		14'h10d9: data = 9'o673;
		14'h10da: data = 9'o372;
		14'h10db: data = 9'o272;
		14'h10dc: data = 9'o172;
		14'h10dd: data = 9'o172;
		14'h10de: data = 9'o272;
		14'h10df: data = 9'o272;
		14'h10e0: data = 9'o272;
		14'h10e1: data = 9'o152;
		14'h10e2: data = 9'o31;
		14'h10e3: data = 9'o41;
		14'h10e4: data = 9'o162;
		14'h10e5: data = 9'o272;
		14'h10e6: data = 9'o272;
		14'h10e7: data = 9'o172;
		14'h10e8: data = 9'o172;
		14'h10e9: data = 9'o272;
		14'h10ea: data = 9'o473;
		14'h10eb: data = 9'o673;
		14'h10ec: data = 9'o773;
		14'h10ed: data = 9'o773;
		14'h10ee: data = 9'o773;
		14'h10ef: data = 9'o773;
		14'h10f0: data = 9'o773;
		14'h10f1: data = 9'o773;
		14'h10f2: data = 9'o363;
		14'h10f3: data = 9'o152;
		14'h10f4: data = 9'o152;
		14'h10f5: data = 9'o152;
		14'h10f6: data = 9'o152;
		14'h10f7: data = 9'o152;
		14'h10f8: data = 9'o152;
		14'h10f9: data = 9'o152;
		14'h10fa: data = 9'o152;
		14'h10fb: data = 9'o152;
		14'h10fc: data = 9'o152;
		14'h10fd: data = 9'o152;
		14'h10fe: data = 9'o152;
		14'h10ff: data = 9'o52;
		14'h1100: data = 9'o52;
		14'h1101: data = 9'o52;
		14'h1102: data = 9'o152;
		14'h1103: data = 9'o152;
		14'h1104: data = 9'o152;
		14'h1105: data = 9'o152;
		14'h1106: data = 9'o142;
		14'h1107: data = 9'o463;
		14'h1108: data = 9'o773;
		14'h1109: data = 9'o773;
		14'h110a: data = 9'o773;
		14'h110b: data = 9'o773;
		14'h110c: data = 9'o773;
		14'h110d: data = 9'o773;
		14'h110e: data = 9'o773;
		14'h110f: data = 9'o473;
		14'h1110: data = 9'o272;
		14'h1111: data = 9'o272;
		14'h1112: data = 9'o172;
		14'h1113: data = 9'o272;
		14'h1114: data = 9'o272;
		14'h1115: data = 9'o162;
		14'h1116: data = 9'o41;
		14'h1117: data = 9'o41;
		14'h1118: data = 9'o152;
		14'h1119: data = 9'o272;
		14'h111a: data = 9'o272;
		14'h111b: data = 9'o172;
		14'h111c: data = 9'o172;
		14'h111d: data = 9'o172;
		14'h111e: data = 9'o172;
		14'h111f: data = 9'o372;
		14'h1120: data = 9'o673;
		14'h1121: data = 9'o773;
		14'h1122: data = 9'o773;
		14'h1123: data = 9'o773;
		14'h1124: data = 9'o773;
		14'h1125: data = 9'o662;
		14'h1126: data = 9'o0;
		14'h1127: data = 9'o0;
		14'h1128: data = 9'o0;
		14'h1129: data = 9'o0;
		14'h112a: data = 9'o0;
		14'h112b: data = 9'o0;
		14'h112c: data = 9'o0;
		14'h112d: data = 9'o0;
		14'h112e: data = 9'o0;
		14'h112f: data = 9'o0;
		14'h1130: data = 9'o0;
		14'h1131: data = 9'o0;
		14'h1132: data = 9'o0;
		14'h1133: data = 9'o0;
		14'h1134: data = 9'o0;
		14'h1135: data = 9'o0;
		14'h1136: data = 9'o0;
		14'h1137: data = 9'o651;
		14'h1138: data = 9'o762;
		14'h1139: data = 9'o773;
		14'h113a: data = 9'o773;
		14'h113b: data = 9'o773;
		14'h113c: data = 9'o773;
		14'h113d: data = 9'o673;
		14'h113e: data = 9'o372;
		14'h113f: data = 9'o272;
		14'h1140: data = 9'o272;
		14'h1141: data = 9'o272;
		14'h1142: data = 9'o272;
		14'h1143: data = 9'o373;
		14'h1144: data = 9'o41;
		14'h1145: data = 9'o20;
		14'h1146: data = 9'o20;
		14'h1147: data = 9'o20;
		14'h1148: data = 9'o31;
		14'h1149: data = 9'o152;
		14'h114a: data = 9'o273;
		14'h114b: data = 9'o172;
		14'h114c: data = 9'o172;
		14'h114d: data = 9'o272;
		14'h114e: data = 9'o372;
		14'h114f: data = 9'o673;
		14'h1150: data = 9'o773;
		14'h1151: data = 9'o773;
		14'h1152: data = 9'o773;
		14'h1153: data = 9'o773;
		14'h1154: data = 9'o773;
		14'h1155: data = 9'o773;
		14'h1156: data = 9'o473;
		14'h1157: data = 9'o152;
		14'h1158: data = 9'o152;
		14'h1159: data = 9'o152;
		14'h115a: data = 9'o152;
		14'h115b: data = 9'o152;
		14'h115c: data = 9'o152;
		14'h115d: data = 9'o152;
		14'h115e: data = 9'o152;
		14'h115f: data = 9'o142;
		14'h1160: data = 9'o142;
		14'h1161: data = 9'o142;
		14'h1162: data = 9'o142;
		14'h1163: data = 9'o152;
		14'h1164: data = 9'o152;
		14'h1165: data = 9'o152;
		14'h1166: data = 9'o152;
		14'h1167: data = 9'o152;
		14'h1168: data = 9'o152;
		14'h1169: data = 9'o252;
		14'h116a: data = 9'o242;
		14'h116b: data = 9'o463;
		14'h116c: data = 9'o773;
		14'h116d: data = 9'o773;
		14'h116e: data = 9'o773;
		14'h116f: data = 9'o773;
		14'h1170: data = 9'o773;
		14'h1171: data = 9'o773;
		14'h1172: data = 9'o673;
		14'h1173: data = 9'o473;
		14'h1174: data = 9'o272;
		14'h1175: data = 9'o272;
		14'h1176: data = 9'o272;
		14'h1177: data = 9'o272;
		14'h1178: data = 9'o262;
		14'h1179: data = 9'o31;
		14'h117a: data = 9'o10;
		14'h117b: data = 9'o10;
		14'h117c: data = 9'o20;
		14'h117d: data = 9'o41;
		14'h117e: data = 9'o272;
		14'h117f: data = 9'o272;
		14'h1180: data = 9'o172;
		14'h1181: data = 9'o172;
		14'h1182: data = 9'o272;
		14'h1183: data = 9'o272;
		14'h1184: data = 9'o673;
		14'h1185: data = 9'o773;
		14'h1186: data = 9'o773;
		14'h1187: data = 9'o773;
		14'h1188: data = 9'o773;
		14'h1189: data = 9'o662;
		14'h118a: data = 9'o0;
		14'h118b: data = 9'o0;
		14'h118c: data = 9'o0;
		14'h118d: data = 9'o0;
		14'h118e: data = 9'o0;
		14'h118f: data = 9'o0;
		14'h1190: data = 9'o0;
		14'h1191: data = 9'o0;
		14'h1192: data = 9'o0;
		14'h1193: data = 9'o0;
		14'h1194: data = 9'o0;
		14'h1195: data = 9'o0;
		14'h1196: data = 9'o0;
		14'h1197: data = 9'o0;
		14'h1198: data = 9'o0;
		14'h1199: data = 9'o0;
		14'h119a: data = 9'o0;
		14'h119b: data = 9'o651;
		14'h119c: data = 9'o762;
		14'h119d: data = 9'o773;
		14'h119e: data = 9'o773;
		14'h119f: data = 9'o773;
		14'h11a0: data = 9'o773;
		14'h11a1: data = 9'o573;
		14'h11a2: data = 9'o272;
		14'h11a3: data = 9'o272;
		14'h11a4: data = 9'o272;
		14'h11a5: data = 9'o272;
		14'h11a6: data = 9'o272;
		14'h11a7: data = 9'o252;
		14'h11a8: data = 9'o20;
		14'h11a9: data = 9'o10;
		14'h11aa: data = 9'o20;
		14'h11ab: data = 9'o10;
		14'h11ac: data = 9'o10;
		14'h11ad: data = 9'o31;
		14'h11ae: data = 9'o272;
		14'h11af: data = 9'o272;
		14'h11b0: data = 9'o172;
		14'h11b1: data = 9'o272;
		14'h11b2: data = 9'o272;
		14'h11b3: data = 9'o573;
		14'h11b4: data = 9'o773;
		14'h11b5: data = 9'o773;
		14'h11b6: data = 9'o773;
		14'h11b7: data = 9'o773;
		14'h11b8: data = 9'o773;
		14'h11b9: data = 9'o773;
		14'h11ba: data = 9'o463;
		14'h11bb: data = 9'o252;
		14'h11bc: data = 9'o152;
		14'h11bd: data = 9'o152;
		14'h11be: data = 9'o152;
		14'h11bf: data = 9'o152;
		14'h11c0: data = 9'o152;
		14'h11c1: data = 9'o142;
		14'h11c2: data = 9'o31;
		14'h11c3: data = 9'o21;
		14'h11c4: data = 9'o21;
		14'h11c5: data = 9'o10;
		14'h11c6: data = 9'o21;
		14'h11c7: data = 9'o31;
		14'h11c8: data = 9'o142;
		14'h11c9: data = 9'o152;
		14'h11ca: data = 9'o152;
		14'h11cb: data = 9'o152;
		14'h11cc: data = 9'o152;
		14'h11cd: data = 9'o242;
		14'h11ce: data = 9'o242;
		14'h11cf: data = 9'o463;
		14'h11d0: data = 9'o773;
		14'h11d1: data = 9'o773;
		14'h11d2: data = 9'o773;
		14'h11d3: data = 9'o773;
		14'h11d4: data = 9'o773;
		14'h11d5: data = 9'o773;
		14'h11d6: data = 9'o673;
		14'h11d7: data = 9'o372;
		14'h11d8: data = 9'o272;
		14'h11d9: data = 9'o172;
		14'h11da: data = 9'o272;
		14'h11db: data = 9'o262;
		14'h11dc: data = 9'o31;
		14'h11dd: data = 9'o10;
		14'h11de: data = 9'o10;
		14'h11df: data = 9'o20;
		14'h11e0: data = 9'o10;
		14'h11e1: data = 9'o20;
		14'h11e2: data = 9'o152;
		14'h11e3: data = 9'o273;
		14'h11e4: data = 9'o172;
		14'h11e5: data = 9'o172;
		14'h11e6: data = 9'o272;
		14'h11e7: data = 9'o272;
		14'h11e8: data = 9'o573;
		14'h11e9: data = 9'o773;
		14'h11ea: data = 9'o773;
		14'h11eb: data = 9'o773;
		14'h11ec: data = 9'o773;
		14'h11ed: data = 9'o662;
		14'h11ee: data = 9'o0;
		14'h11ef: data = 9'o0;
		14'h11f0: data = 9'o0;
		14'h11f1: data = 9'o0;
		14'h11f2: data = 9'o0;
		14'h11f3: data = 9'o0;
		14'h11f4: data = 9'o0;
		14'h11f5: data = 9'o0;
		14'h11f6: data = 9'o0;
		14'h11f7: data = 9'o0;
		14'h11f8: data = 9'o0;
		14'h11f9: data = 9'o0;
		14'h11fa: data = 9'o0;
		14'h11fb: data = 9'o0;
		14'h11fc: data = 9'o0;
		14'h11fd: data = 9'o0;
		14'h11fe: data = 9'o0;
		14'h11ff: data = 9'o651;
		14'h1200: data = 9'o762;
		14'h1201: data = 9'o773;
		14'h1202: data = 9'o773;
		14'h1203: data = 9'o773;
		14'h1204: data = 9'o773;
		14'h1205: data = 9'o573;
		14'h1206: data = 9'o272;
		14'h1207: data = 9'o172;
		14'h1208: data = 9'o172;
		14'h1209: data = 9'o273;
		14'h120a: data = 9'o272;
		14'h120b: data = 9'o31;
		14'h120c: data = 9'o10;
		14'h120d: data = 9'o10;
		14'h120e: data = 9'o10;
		14'h120f: data = 9'o10;
		14'h1210: data = 9'o10;
		14'h1211: data = 9'o20;
		14'h1212: data = 9'o152;
		14'h1213: data = 9'o273;
		14'h1214: data = 9'o272;
		14'h1215: data = 9'o172;
		14'h1216: data = 9'o272;
		14'h1217: data = 9'o473;
		14'h1218: data = 9'o773;
		14'h1219: data = 9'o773;
		14'h121a: data = 9'o773;
		14'h121b: data = 9'o773;
		14'h121c: data = 9'o773;
		14'h121d: data = 9'o773;
		14'h121e: data = 9'o673;
		14'h121f: data = 9'o573;
		14'h1220: data = 9'o573;
		14'h1221: data = 9'o373;
		14'h1222: data = 9'o152;
		14'h1223: data = 9'o152;
		14'h1224: data = 9'o152;
		14'h1225: data = 9'o31;
		14'h1226: data = 9'o21;
		14'h1227: data = 9'o10;
		14'h1228: data = 9'o10;
		14'h1229: data = 9'o10;
		14'h122a: data = 9'o10;
		14'h122b: data = 9'o21;
		14'h122c: data = 9'o31;
		14'h122d: data = 9'o152;
		14'h122e: data = 9'o152;
		14'h122f: data = 9'o152;
		14'h1230: data = 9'o363;
		14'h1231: data = 9'o573;
		14'h1232: data = 9'o573;
		14'h1233: data = 9'o673;
		14'h1234: data = 9'o773;
		14'h1235: data = 9'o773;
		14'h1236: data = 9'o773;
		14'h1237: data = 9'o773;
		14'h1238: data = 9'o773;
		14'h1239: data = 9'o773;
		14'h123a: data = 9'o573;
		14'h123b: data = 9'o272;
		14'h123c: data = 9'o272;
		14'h123d: data = 9'o272;
		14'h123e: data = 9'o172;
		14'h123f: data = 9'o162;
		14'h1240: data = 9'o20;
		14'h1241: data = 9'o10;
		14'h1242: data = 9'o10;
		14'h1243: data = 9'o10;
		14'h1244: data = 9'o10;
		14'h1245: data = 9'o20;
		14'h1246: data = 9'o31;
		14'h1247: data = 9'o272;
		14'h1248: data = 9'o272;
		14'h1249: data = 9'o172;
		14'h124a: data = 9'o272;
		14'h124b: data = 9'o272;
		14'h124c: data = 9'o573;
		14'h124d: data = 9'o773;
		14'h124e: data = 9'o773;
		14'h124f: data = 9'o773;
		14'h1250: data = 9'o773;
		14'h1251: data = 9'o662;
		14'h1252: data = 9'o0;
		14'h1253: data = 9'o0;
		14'h1254: data = 9'o0;
		14'h1255: data = 9'o0;
		14'h1256: data = 9'o0;
		14'h1257: data = 9'o0;
		14'h1258: data = 9'o0;
		14'h1259: data = 9'o0;
		14'h125a: data = 9'o0;
		14'h125b: data = 9'o0;
		14'h125c: data = 9'o0;
		14'h125d: data = 9'o0;
		14'h125e: data = 9'o0;
		14'h125f: data = 9'o0;
		14'h1260: data = 9'o0;
		14'h1261: data = 9'o0;
		14'h1262: data = 9'o0;
		14'h1263: data = 9'o651;
		14'h1264: data = 9'o762;
		14'h1265: data = 9'o773;
		14'h1266: data = 9'o773;
		14'h1267: data = 9'o773;
		14'h1268: data = 9'o673;
		14'h1269: data = 9'o473;
		14'h126a: data = 9'o272;
		14'h126b: data = 9'o172;
		14'h126c: data = 9'o172;
		14'h126d: data = 9'o273;
		14'h126e: data = 9'o262;
		14'h126f: data = 9'o20;
		14'h1270: data = 9'o10;
		14'h1271: data = 9'o10;
		14'h1272: data = 9'o10;
		14'h1273: data = 9'o11;
		14'h1274: data = 9'o10;
		14'h1275: data = 9'o10;
		14'h1276: data = 9'o31;
		14'h1277: data = 9'o272;
		14'h1278: data = 9'o273;
		14'h1279: data = 9'o272;
		14'h127a: data = 9'o272;
		14'h127b: data = 9'o473;
		14'h127c: data = 9'o773;
		14'h127d: data = 9'o773;
		14'h127e: data = 9'o773;
		14'h127f: data = 9'o773;
		14'h1280: data = 9'o773;
		14'h1281: data = 9'o773;
		14'h1282: data = 9'o773;
		14'h1283: data = 9'o773;
		14'h1284: data = 9'o773;
		14'h1285: data = 9'o573;
		14'h1286: data = 9'o152;
		14'h1287: data = 9'o152;
		14'h1288: data = 9'o142;
		14'h1289: data = 9'o21;
		14'h128a: data = 9'o10;
		14'h128b: data = 9'o10;
		14'h128c: data = 9'o11;
		14'h128d: data = 9'o10;
		14'h128e: data = 9'o10;
		14'h128f: data = 9'o10;
		14'h1290: data = 9'o21;
		14'h1291: data = 9'o142;
		14'h1292: data = 9'o152;
		14'h1293: data = 9'o152;
		14'h1294: data = 9'o473;
		14'h1295: data = 9'o773;
		14'h1296: data = 9'o773;
		14'h1297: data = 9'o773;
		14'h1298: data = 9'o773;
		14'h1299: data = 9'o773;
		14'h129a: data = 9'o773;
		14'h129b: data = 9'o773;
		14'h129c: data = 9'o773;
		14'h129d: data = 9'o773;
		14'h129e: data = 9'o473;
		14'h129f: data = 9'o272;
		14'h12a0: data = 9'o272;
		14'h12a1: data = 9'o272;
		14'h12a2: data = 9'o272;
		14'h12a3: data = 9'o41;
		14'h12a4: data = 9'o10;
		14'h12a5: data = 9'o10;
		14'h12a6: data = 9'o10;
		14'h12a7: data = 9'o10;
		14'h12a8: data = 9'o10;
		14'h12a9: data = 9'o10;
		14'h12aa: data = 9'o20;
		14'h12ab: data = 9'o152;
		14'h12ac: data = 9'o273;
		14'h12ad: data = 9'o172;
		14'h12ae: data = 9'o272;
		14'h12af: data = 9'o272;
		14'h12b0: data = 9'o473;
		14'h12b1: data = 9'o773;
		14'h12b2: data = 9'o773;
		14'h12b3: data = 9'o773;
		14'h12b4: data = 9'o773;
		14'h12b5: data = 9'o662;
		14'h12b6: data = 9'o0;
		14'h12b7: data = 9'o0;
		14'h12b8: data = 9'o0;
		14'h12b9: data = 9'o0;
		14'h12ba: data = 9'o0;
		14'h12bb: data = 9'o0;
		14'h12bc: data = 9'o0;
		14'h12bd: data = 9'o0;
		14'h12be: data = 9'o0;
		14'h12bf: data = 9'o0;
		14'h12c0: data = 9'o0;
		14'h12c1: data = 9'o0;
		14'h12c2: data = 9'o0;
		14'h12c3: data = 9'o0;
		14'h12c4: data = 9'o0;
		14'h12c5: data = 9'o0;
		14'h12c6: data = 9'o0;
		14'h12c7: data = 9'o651;
		14'h12c8: data = 9'o762;
		14'h12c9: data = 9'o773;
		14'h12ca: data = 9'o773;
		14'h12cb: data = 9'o773;
		14'h12cc: data = 9'o673;
		14'h12cd: data = 9'o473;
		14'h12ce: data = 9'o272;
		14'h12cf: data = 9'o172;
		14'h12d0: data = 9'o172;
		14'h12d1: data = 9'o273;
		14'h12d2: data = 9'o41;
		14'h12d3: data = 9'o10;
		14'h12d4: data = 9'o10;
		14'h12d5: data = 9'o10;
		14'h12d6: data = 9'o10;
		14'h12d7: data = 9'o10;
		14'h12d8: data = 9'o10;
		14'h12d9: data = 9'o10;
		14'h12da: data = 9'o20;
		14'h12db: data = 9'o262;
		14'h12dc: data = 9'o272;
		14'h12dd: data = 9'o272;
		14'h12de: data = 9'o272;
		14'h12df: data = 9'o473;
		14'h12e0: data = 9'o773;
		14'h12e1: data = 9'o773;
		14'h12e2: data = 9'o773;
		14'h12e3: data = 9'o773;
		14'h12e4: data = 9'o773;
		14'h12e5: data = 9'o773;
		14'h12e6: data = 9'o773;
		14'h12e7: data = 9'o773;
		14'h12e8: data = 9'o773;
		14'h12e9: data = 9'o573;
		14'h12ea: data = 9'o252;
		14'h12eb: data = 9'o152;
		14'h12ec: data = 9'o142;
		14'h12ed: data = 9'o21;
		14'h12ee: data = 9'o11;
		14'h12ef: data = 9'o10;
		14'h12f0: data = 9'o10;
		14'h12f1: data = 9'o10;
		14'h12f2: data = 9'o10;
		14'h12f3: data = 9'o10;
		14'h12f4: data = 9'o10;
		14'h12f5: data = 9'o42;
		14'h12f6: data = 9'o152;
		14'h12f7: data = 9'o152;
		14'h12f8: data = 9'o563;
		14'h12f9: data = 9'o773;
		14'h12fa: data = 9'o773;
		14'h12fb: data = 9'o773;
		14'h12fc: data = 9'o773;
		14'h12fd: data = 9'o773;
		14'h12fe: data = 9'o773;
		14'h12ff: data = 9'o773;
		14'h1300: data = 9'o773;
		14'h1301: data = 9'o773;
		14'h1302: data = 9'o473;
		14'h1303: data = 9'o272;
		14'h1304: data = 9'o272;
		14'h1305: data = 9'o272;
		14'h1306: data = 9'o272;
		14'h1307: data = 9'o20;
		14'h1308: data = 9'o20;
		14'h1309: data = 9'o10;
		14'h130a: data = 9'o10;
		14'h130b: data = 9'o10;
		14'h130c: data = 9'o11;
		14'h130d: data = 9'o10;
		14'h130e: data = 9'o20;
		14'h130f: data = 9'o41;
		14'h1310: data = 9'o272;
		14'h1311: data = 9'o172;
		14'h1312: data = 9'o272;
		14'h1313: data = 9'o272;
		14'h1314: data = 9'o473;
		14'h1315: data = 9'o673;
		14'h1316: data = 9'o773;
		14'h1317: data = 9'o773;
		14'h1318: data = 9'o773;
		14'h1319: data = 9'o662;
		14'h131a: data = 9'o0;
		14'h131b: data = 9'o0;
		14'h131c: data = 9'o0;
		14'h131d: data = 9'o0;
		14'h131e: data = 9'o0;
		14'h131f: data = 9'o0;
		14'h1320: data = 9'o0;
		14'h1321: data = 9'o0;
		14'h1322: data = 9'o0;
		14'h1323: data = 9'o0;
		14'h1324: data = 9'o0;
		14'h1325: data = 9'o0;
		14'h1326: data = 9'o0;
		14'h1327: data = 9'o0;
		14'h1328: data = 9'o0;
		14'h1329: data = 9'o0;
		14'h132a: data = 9'o0;
		14'h132b: data = 9'o651;
		14'h132c: data = 9'o762;
		14'h132d: data = 9'o773;
		14'h132e: data = 9'o773;
		14'h132f: data = 9'o773;
		14'h1330: data = 9'o673;
		14'h1331: data = 9'o373;
		14'h1332: data = 9'o272;
		14'h1333: data = 9'o172;
		14'h1334: data = 9'o172;
		14'h1335: data = 9'o273;
		14'h1336: data = 9'o31;
		14'h1337: data = 9'o10;
		14'h1338: data = 9'o10;
		14'h1339: data = 9'o10;
		14'h133a: data = 9'o11;
		14'h133b: data = 9'o10;
		14'h133c: data = 9'o10;
		14'h133d: data = 9'o10;
		14'h133e: data = 9'o20;
		14'h133f: data = 9'o152;
		14'h1340: data = 9'o273;
		14'h1341: data = 9'o172;
		14'h1342: data = 9'o272;
		14'h1343: data = 9'o372;
		14'h1344: data = 9'o673;
		14'h1345: data = 9'o773;
		14'h1346: data = 9'o773;
		14'h1347: data = 9'o773;
		14'h1348: data = 9'o773;
		14'h1349: data = 9'o773;
		14'h134a: data = 9'o773;
		14'h134b: data = 9'o773;
		14'h134c: data = 9'o773;
		14'h134d: data = 9'o573;
		14'h134e: data = 9'o142;
		14'h134f: data = 9'o152;
		14'h1350: data = 9'o142;
		14'h1351: data = 9'o11;
		14'h1352: data = 9'o11;
		14'h1353: data = 9'o10;
		14'h1354: data = 9'o10;
		14'h1355: data = 9'o10;
		14'h1356: data = 9'o11;
		14'h1357: data = 9'o10;
		14'h1358: data = 9'o10;
		14'h1359: data = 9'o42;
		14'h135a: data = 9'o52;
		14'h135b: data = 9'o152;
		14'h135c: data = 9'o463;
		14'h135d: data = 9'o773;
		14'h135e: data = 9'o773;
		14'h135f: data = 9'o773;
		14'h1360: data = 9'o773;
		14'h1361: data = 9'o773;
		14'h1362: data = 9'o773;
		14'h1363: data = 9'o773;
		14'h1364: data = 9'o773;
		14'h1365: data = 9'o673;
		14'h1366: data = 9'o373;
		14'h1367: data = 9'o272;
		14'h1368: data = 9'o272;
		14'h1369: data = 9'o272;
		14'h136a: data = 9'o162;
		14'h136b: data = 9'o20;
		14'h136c: data = 9'o10;
		14'h136d: data = 9'o11;
		14'h136e: data = 9'o10;
		14'h136f: data = 9'o10;
		14'h1370: data = 9'o10;
		14'h1371: data = 9'o10;
		14'h1372: data = 9'o10;
		14'h1373: data = 9'o20;
		14'h1374: data = 9'o272;
		14'h1375: data = 9'o172;
		14'h1376: data = 9'o172;
		14'h1377: data = 9'o272;
		14'h1378: data = 9'o373;
		14'h1379: data = 9'o673;
		14'h137a: data = 9'o773;
		14'h137b: data = 9'o773;
		14'h137c: data = 9'o773;
		14'h137d: data = 9'o662;
		14'h137e: data = 9'o0;
		14'h137f: data = 9'o0;
		14'h1380: data = 9'o0;
		14'h1381: data = 9'o0;
		14'h1382: data = 9'o0;
		14'h1383: data = 9'o0;
		14'h1384: data = 9'o0;
		14'h1385: data = 9'o0;
		14'h1386: data = 9'o0;
		14'h1387: data = 9'o0;
		14'h1388: data = 9'o0;
		14'h1389: data = 9'o0;
		14'h138a: data = 9'o0;
		14'h138b: data = 9'o0;
		14'h138c: data = 9'o0;
		14'h138d: data = 9'o0;
		14'h138e: data = 9'o0;
		14'h138f: data = 9'o651;
		14'h1390: data = 9'o662;
		14'h1391: data = 9'o773;
		14'h1392: data = 9'o773;
		14'h1393: data = 9'o773;
		14'h1394: data = 9'o673;
		14'h1395: data = 9'o372;
		14'h1396: data = 9'o272;
		14'h1397: data = 9'o172;
		14'h1398: data = 9'o172;
		14'h1399: data = 9'o162;
		14'h139a: data = 9'o20;
		14'h139b: data = 9'o10;
		14'h139c: data = 9'o10;
		14'h139d: data = 9'o10;
		14'h139e: data = 9'o10;
		14'h139f: data = 9'o10;
		14'h13a0: data = 9'o10;
		14'h13a1: data = 9'o10;
		14'h13a2: data = 9'o10;
		14'h13a3: data = 9'o41;
		14'h13a4: data = 9'o272;
		14'h13a5: data = 9'o172;
		14'h13a6: data = 9'o272;
		14'h13a7: data = 9'o373;
		14'h13a8: data = 9'o673;
		14'h13a9: data = 9'o673;
		14'h13aa: data = 9'o773;
		14'h13ab: data = 9'o773;
		14'h13ac: data = 9'o773;
		14'h13ad: data = 9'o773;
		14'h13ae: data = 9'o773;
		14'h13af: data = 9'o773;
		14'h13b0: data = 9'o673;
		14'h13b1: data = 9'o573;
		14'h13b2: data = 9'o152;
		14'h13b3: data = 9'o152;
		14'h13b4: data = 9'o142;
		14'h13b5: data = 9'o21;
		14'h13b6: data = 9'o11;
		14'h13b7: data = 9'o10;
		14'h13b8: data = 9'o11;
		14'h13b9: data = 9'o10;
		14'h13ba: data = 9'o10;
		14'h13bb: data = 9'o10;
		14'h13bc: data = 9'o21;
		14'h13bd: data = 9'o42;
		14'h13be: data = 9'o152;
		14'h13bf: data = 9'o152;
		14'h13c0: data = 9'o473;
		14'h13c1: data = 9'o673;
		14'h13c2: data = 9'o773;
		14'h13c3: data = 9'o773;
		14'h13c4: data = 9'o773;
		14'h13c5: data = 9'o773;
		14'h13c6: data = 9'o773;
		14'h13c7: data = 9'o773;
		14'h13c8: data = 9'o773;
		14'h13c9: data = 9'o673;
		14'h13ca: data = 9'o373;
		14'h13cb: data = 9'o272;
		14'h13cc: data = 9'o172;
		14'h13cd: data = 9'o272;
		14'h13ce: data = 9'o41;
		14'h13cf: data = 9'o20;
		14'h13d0: data = 9'o10;
		14'h13d1: data = 9'o10;
		14'h13d2: data = 9'o10;
		14'h13d3: data = 9'o10;
		14'h13d4: data = 9'o10;
		14'h13d5: data = 9'o10;
		14'h13d6: data = 9'o10;
		14'h13d7: data = 9'o20;
		14'h13d8: data = 9'o162;
		14'h13d9: data = 9'o272;
		14'h13da: data = 9'o172;
		14'h13db: data = 9'o272;
		14'h13dc: data = 9'o372;
		14'h13dd: data = 9'o673;
		14'h13de: data = 9'o773;
		14'h13df: data = 9'o773;
		14'h13e0: data = 9'o773;
		14'h13e1: data = 9'o662;
		14'h13e2: data = 9'o0;
		14'h13e3: data = 9'o0;
		14'h13e4: data = 9'o0;
		14'h13e5: data = 9'o0;
		14'h13e6: data = 9'o0;
		14'h13e7: data = 9'o0;
		14'h13e8: data = 9'o0;
		14'h13e9: data = 9'o0;
		14'h13ea: data = 9'o0;
		14'h13eb: data = 9'o0;
		14'h13ec: data = 9'o0;
		14'h13ed: data = 9'o0;
		14'h13ee: data = 9'o0;
		14'h13ef: data = 9'o0;
		14'h13f0: data = 9'o0;
		14'h13f1: data = 9'o0;
		14'h13f2: data = 9'o0;
		14'h13f3: data = 9'o651;
		14'h13f4: data = 9'o662;
		14'h13f5: data = 9'o773;
		14'h13f6: data = 9'o773;
		14'h13f7: data = 9'o773;
		14'h13f8: data = 9'o673;
		14'h13f9: data = 9'o372;
		14'h13fa: data = 9'o272;
		14'h13fb: data = 9'o272;
		14'h13fc: data = 9'o273;
		14'h13fd: data = 9'o152;
		14'h13fe: data = 9'o20;
		14'h13ff: data = 9'o10;
		14'h1400: data = 9'o10;
		14'h1401: data = 9'o10;
		14'h1402: data = 9'o10;
		14'h1403: data = 9'o10;
		14'h1404: data = 9'o10;
		14'h1405: data = 9'o10;
		14'h1406: data = 9'o20;
		14'h1407: data = 9'o31;
		14'h1408: data = 9'o272;
		14'h1409: data = 9'o172;
		14'h140a: data = 9'o172;
		14'h140b: data = 9'o272;
		14'h140c: data = 9'o473;
		14'h140d: data = 9'o573;
		14'h140e: data = 9'o573;
		14'h140f: data = 9'o773;
		14'h1410: data = 9'o773;
		14'h1411: data = 9'o773;
		14'h1412: data = 9'o673;
		14'h1413: data = 9'o473;
		14'h1414: data = 9'o473;
		14'h1415: data = 9'o373;
		14'h1416: data = 9'o152;
		14'h1417: data = 9'o152;
		14'h1418: data = 9'o142;
		14'h1419: data = 9'o31;
		14'h141a: data = 9'o11;
		14'h141b: data = 9'o11;
		14'h141c: data = 9'o11;
		14'h141d: data = 9'o10;
		14'h141e: data = 9'o10;
		14'h141f: data = 9'o21;
		14'h1420: data = 9'o31;
		14'h1421: data = 9'o152;
		14'h1422: data = 9'o152;
		14'h1423: data = 9'o152;
		14'h1424: data = 9'o373;
		14'h1425: data = 9'o473;
		14'h1426: data = 9'o573;
		14'h1427: data = 9'o673;
		14'h1428: data = 9'o773;
		14'h1429: data = 9'o773;
		14'h142a: data = 9'o773;
		14'h142b: data = 9'o673;
		14'h142c: data = 9'o573;
		14'h142d: data = 9'o473;
		14'h142e: data = 9'o272;
		14'h142f: data = 9'o172;
		14'h1430: data = 9'o172;
		14'h1431: data = 9'o272;
		14'h1432: data = 9'o31;
		14'h1433: data = 9'o10;
		14'h1434: data = 9'o10;
		14'h1435: data = 9'o10;
		14'h1436: data = 9'o10;
		14'h1437: data = 9'o11;
		14'h1438: data = 9'o10;
		14'h1439: data = 9'o10;
		14'h143a: data = 9'o10;
		14'h143b: data = 9'o10;
		14'h143c: data = 9'o51;
		14'h143d: data = 9'o272;
		14'h143e: data = 9'o172;
		14'h143f: data = 9'o272;
		14'h1440: data = 9'o372;
		14'h1441: data = 9'o673;
		14'h1442: data = 9'o773;
		14'h1443: data = 9'o773;
		14'h1444: data = 9'o773;
		14'h1445: data = 9'o762;
		14'h1446: data = 9'o0;
		14'h1447: data = 9'o0;
		14'h1448: data = 9'o0;
		14'h1449: data = 9'o0;
		14'h144a: data = 9'o0;
		14'h144b: data = 9'o0;
		14'h144c: data = 9'o0;
		14'h144d: data = 9'o0;
		14'h144e: data = 9'o0;
		14'h144f: data = 9'o0;
		14'h1450: data = 9'o0;
		14'h1451: data = 9'o0;
		14'h1452: data = 9'o0;
		14'h1453: data = 9'o0;
		14'h1454: data = 9'o0;
		14'h1455: data = 9'o0;
		14'h1456: data = 9'o0;
		14'h1457: data = 9'o551;
		14'h1458: data = 9'o662;
		14'h1459: data = 9'o773;
		14'h145a: data = 9'o773;
		14'h145b: data = 9'o773;
		14'h145c: data = 9'o573;
		14'h145d: data = 9'o372;
		14'h145e: data = 9'o272;
		14'h145f: data = 9'o272;
		14'h1460: data = 9'o272;
		14'h1461: data = 9'o41;
		14'h1462: data = 9'o20;
		14'h1463: data = 9'o10;
		14'h1464: data = 9'o10;
		14'h1465: data = 9'o10;
		14'h1466: data = 9'o10;
		14'h1467: data = 9'o10;
		14'h1468: data = 9'o10;
		14'h1469: data = 9'o10;
		14'h146a: data = 9'o10;
		14'h146b: data = 9'o20;
		14'h146c: data = 9'o162;
		14'h146d: data = 9'o172;
		14'h146e: data = 9'o172;
		14'h146f: data = 9'o172;
		14'h1470: data = 9'o272;
		14'h1471: data = 9'o372;
		14'h1472: data = 9'o473;
		14'h1473: data = 9'o673;
		14'h1474: data = 9'o773;
		14'h1475: data = 9'o773;
		14'h1476: data = 9'o473;
		14'h1477: data = 9'o372;
		14'h1478: data = 9'o273;
		14'h1479: data = 9'o263;
		14'h147a: data = 9'o52;
		14'h147b: data = 9'o152;
		14'h147c: data = 9'o152;
		14'h147d: data = 9'o142;
		14'h147e: data = 9'o21;
		14'h147f: data = 9'o21;
		14'h1480: data = 9'o11;
		14'h1481: data = 9'o10;
		14'h1482: data = 9'o21;
		14'h1483: data = 9'o31;
		14'h1484: data = 9'o142;
		14'h1485: data = 9'o152;
		14'h1486: data = 9'o152;
		14'h1487: data = 9'o152;
		14'h1488: data = 9'o262;
		14'h1489: data = 9'o273;
		14'h148a: data = 9'o372;
		14'h148b: data = 9'o573;
		14'h148c: data = 9'o773;
		14'h148d: data = 9'o773;
		14'h148e: data = 9'o673;
		14'h148f: data = 9'o473;
		14'h1490: data = 9'o372;
		14'h1491: data = 9'o272;
		14'h1492: data = 9'o172;
		14'h1493: data = 9'o172;
		14'h1494: data = 9'o172;
		14'h1495: data = 9'o272;
		14'h1496: data = 9'o20;
		14'h1497: data = 9'o10;
		14'h1498: data = 9'o10;
		14'h1499: data = 9'o10;
		14'h149a: data = 9'o10;
		14'h149b: data = 9'o10;
		14'h149c: data = 9'o10;
		14'h149d: data = 9'o10;
		14'h149e: data = 9'o10;
		14'h149f: data = 9'o10;
		14'h14a0: data = 9'o41;
		14'h14a1: data = 9'o272;
		14'h14a2: data = 9'o272;
		14'h14a3: data = 9'o272;
		14'h14a4: data = 9'o372;
		14'h14a5: data = 9'o573;
		14'h14a6: data = 9'o773;
		14'h14a7: data = 9'o773;
		14'h14a8: data = 9'o773;
		14'h14a9: data = 9'o762;
		14'h14aa: data = 9'o0;
		14'h14ab: data = 9'o0;
		14'h14ac: data = 9'o0;
		14'h14ad: data = 9'o0;
		14'h14ae: data = 9'o0;
		14'h14af: data = 9'o0;
		14'h14b0: data = 9'o0;
		14'h14b1: data = 9'o0;
		14'h14b2: data = 9'o0;
		14'h14b3: data = 9'o0;
		14'h14b4: data = 9'o0;
		14'h14b5: data = 9'o0;
		14'h14b6: data = 9'o0;
		14'h14b7: data = 9'o0;
		14'h14b8: data = 9'o0;
		14'h14b9: data = 9'o0;
		14'h14ba: data = 9'o0;
		14'h14bb: data = 9'o651;
		14'h14bc: data = 9'o662;
		14'h14bd: data = 9'o773;
		14'h14be: data = 9'o773;
		14'h14bf: data = 9'o773;
		14'h14c0: data = 9'o573;
		14'h14c1: data = 9'o372;
		14'h14c2: data = 9'o272;
		14'h14c3: data = 9'o272;
		14'h14c4: data = 9'o272;
		14'h14c5: data = 9'o41;
		14'h14c6: data = 9'o20;
		14'h14c7: data = 9'o10;
		14'h14c8: data = 9'o20;
		14'h14c9: data = 9'o20;
		14'h14ca: data = 9'o20;
		14'h14cb: data = 9'o20;
		14'h14cc: data = 9'o10;
		14'h14cd: data = 9'o10;
		14'h14ce: data = 9'o10;
		14'h14cf: data = 9'o20;
		14'h14d0: data = 9'o152;
		14'h14d1: data = 9'o272;
		14'h14d2: data = 9'o272;
		14'h14d3: data = 9'o272;
		14'h14d4: data = 9'o272;
		14'h14d5: data = 9'o272;
		14'h14d6: data = 9'o473;
		14'h14d7: data = 9'o673;
		14'h14d8: data = 9'o773;
		14'h14d9: data = 9'o773;
		14'h14da: data = 9'o473;
		14'h14db: data = 9'o272;
		14'h14dc: data = 9'o272;
		14'h14dd: data = 9'o162;
		14'h14de: data = 9'o52;
		14'h14df: data = 9'o152;
		14'h14e0: data = 9'o152;
		14'h14e1: data = 9'o152;
		14'h14e2: data = 9'o152;
		14'h14e3: data = 9'o142;
		14'h14e4: data = 9'o142;
		14'h14e5: data = 9'o142;
		14'h14e6: data = 9'o142;
		14'h14e7: data = 9'o152;
		14'h14e8: data = 9'o152;
		14'h14e9: data = 9'o152;
		14'h14ea: data = 9'o152;
		14'h14eb: data = 9'o152;
		14'h14ec: data = 9'o162;
		14'h14ed: data = 9'o272;
		14'h14ee: data = 9'o272;
		14'h14ef: data = 9'o473;
		14'h14f0: data = 9'o673;
		14'h14f1: data = 9'o773;
		14'h14f2: data = 9'o673;
		14'h14f3: data = 9'o473;
		14'h14f4: data = 9'o272;
		14'h14f5: data = 9'o272;
		14'h14f6: data = 9'o272;
		14'h14f7: data = 9'o272;
		14'h14f8: data = 9'o172;
		14'h14f9: data = 9'o162;
		14'h14fa: data = 9'o20;
		14'h14fb: data = 9'o10;
		14'h14fc: data = 9'o10;
		14'h14fd: data = 9'o10;
		14'h14fe: data = 9'o10;
		14'h14ff: data = 9'o20;
		14'h1500: data = 9'o10;
		14'h1501: data = 9'o10;
		14'h1502: data = 9'o10;
		14'h1503: data = 9'o10;
		14'h1504: data = 9'o31;
		14'h1505: data = 9'o272;
		14'h1506: data = 9'o272;
		14'h1507: data = 9'o272;
		14'h1508: data = 9'o272;
		14'h1509: data = 9'o573;
		14'h150a: data = 9'o773;
		14'h150b: data = 9'o773;
		14'h150c: data = 9'o773;
		14'h150d: data = 9'o762;
		14'h150e: data = 9'o0;
		14'h150f: data = 9'o0;
		14'h1510: data = 9'o0;
		14'h1511: data = 9'o0;
		14'h1512: data = 9'o0;
		14'h1513: data = 9'o0;
		14'h1514: data = 9'o0;
		14'h1515: data = 9'o0;
		14'h1516: data = 9'o0;
		14'h1517: data = 9'o0;
		14'h1518: data = 9'o0;
		14'h1519: data = 9'o0;
		14'h151a: data = 9'o0;
		14'h151b: data = 9'o0;
		14'h151c: data = 9'o0;
		14'h151d: data = 9'o0;
		14'h151e: data = 9'o0;
		14'h151f: data = 9'o651;
		14'h1520: data = 9'o662;
		14'h1521: data = 9'o773;
		14'h1522: data = 9'o773;
		14'h1523: data = 9'o773;
		14'h1524: data = 9'o573;
		14'h1525: data = 9'o372;
		14'h1526: data = 9'o272;
		14'h1527: data = 9'o172;
		14'h1528: data = 9'o172;
		14'h1529: data = 9'o41;
		14'h152a: data = 9'o41;
		14'h152b: data = 9'o31;
		14'h152c: data = 9'o31;
		14'h152d: data = 9'o41;
		14'h152e: data = 9'o31;
		14'h152f: data = 9'o31;
		14'h1530: data = 9'o31;
		14'h1531: data = 9'o131;
		14'h1532: data = 9'o131;
		14'h1533: data = 9'o141;
		14'h1534: data = 9'o162;
		14'h1535: data = 9'o272;
		14'h1536: data = 9'o172;
		14'h1537: data = 9'o272;
		14'h1538: data = 9'o272;
		14'h1539: data = 9'o272;
		14'h153a: data = 9'o373;
		14'h153b: data = 9'o573;
		14'h153c: data = 9'o673;
		14'h153d: data = 9'o673;
		14'h153e: data = 9'o373;
		14'h153f: data = 9'o272;
		14'h1540: data = 9'o273;
		14'h1541: data = 9'o173;
		14'h1542: data = 9'o52;
		14'h1543: data = 9'o152;
		14'h1544: data = 9'o52;
		14'h1545: data = 9'o152;
		14'h1546: data = 9'o152;
		14'h1547: data = 9'o152;
		14'h1548: data = 9'o152;
		14'h1549: data = 9'o152;
		14'h154a: data = 9'o152;
		14'h154b: data = 9'o152;
		14'h154c: data = 9'o152;
		14'h154d: data = 9'o52;
		14'h154e: data = 9'o152;
		14'h154f: data = 9'o152;
		14'h1550: data = 9'o162;
		14'h1551: data = 9'o272;
		14'h1552: data = 9'o272;
		14'h1553: data = 9'o373;
		14'h1554: data = 9'o573;
		14'h1555: data = 9'o673;
		14'h1556: data = 9'o573;
		14'h1557: data = 9'o373;
		14'h1558: data = 9'o273;
		14'h1559: data = 9'o272;
		14'h155a: data = 9'o272;
		14'h155b: data = 9'o172;
		14'h155c: data = 9'o172;
		14'h155d: data = 9'o162;
		14'h155e: data = 9'o41;
		14'h155f: data = 9'o31;
		14'h1560: data = 9'o31;
		14'h1561: data = 9'o31;
		14'h1562: data = 9'o31;
		14'h1563: data = 9'o31;
		14'h1564: data = 9'o31;
		14'h1565: data = 9'o31;
		14'h1566: data = 9'o31;
		14'h1567: data = 9'o41;
		14'h1568: data = 9'o41;
		14'h1569: data = 9'o272;
		14'h156a: data = 9'o172;
		14'h156b: data = 9'o272;
		14'h156c: data = 9'o272;
		14'h156d: data = 9'o473;
		14'h156e: data = 9'o773;
		14'h156f: data = 9'o773;
		14'h1570: data = 9'o773;
		14'h1571: data = 9'o762;
		14'h1572: data = 9'o0;
		14'h1573: data = 9'o0;
		14'h1574: data = 9'o0;
		14'h1575: data = 9'o0;
		14'h1576: data = 9'o0;
		14'h1577: data = 9'o0;
		14'h1578: data = 9'o0;
		14'h1579: data = 9'o0;
		14'h157a: data = 9'o0;
		14'h157b: data = 9'o0;
		14'h157c: data = 9'o0;
		14'h157d: data = 9'o0;
		14'h157e: data = 9'o0;
		14'h157f: data = 9'o0;
		14'h1580: data = 9'o0;
		14'h1581: data = 9'o0;
		14'h1582: data = 9'o0;
		14'h1583: data = 9'o651;
		14'h1584: data = 9'o762;
		14'h1585: data = 9'o773;
		14'h1586: data = 9'o773;
		14'h1587: data = 9'o673;
		14'h1588: data = 9'o473;
		14'h1589: data = 9'o272;
		14'h158a: data = 9'o272;
		14'h158b: data = 9'o172;
		14'h158c: data = 9'o173;
		14'h158d: data = 9'o172;
		14'h158e: data = 9'o273;
		14'h158f: data = 9'o272;
		14'h1590: data = 9'o273;
		14'h1591: data = 9'o273;
		14'h1592: data = 9'o273;
		14'h1593: data = 9'o273;
		14'h1594: data = 9'o272;
		14'h1595: data = 9'o272;
		14'h1596: data = 9'o272;
		14'h1597: data = 9'o272;
		14'h1598: data = 9'o172;
		14'h1599: data = 9'o172;
		14'h159a: data = 9'o172;
		14'h159b: data = 9'o272;
		14'h159c: data = 9'o272;
		14'h159d: data = 9'o272;
		14'h159e: data = 9'o272;
		14'h159f: data = 9'o273;
		14'h15a0: data = 9'o373;
		14'h15a1: data = 9'o373;
		14'h15a2: data = 9'o272;
		14'h15a3: data = 9'o272;
		14'h15a4: data = 9'o273;
		14'h15a5: data = 9'o173;
		14'h15a6: data = 9'o152;
		14'h15a7: data = 9'o152;
		14'h15a8: data = 9'o52;
		14'h15a9: data = 9'o152;
		14'h15aa: data = 9'o52;
		14'h15ab: data = 9'o152;
		14'h15ac: data = 9'o152;
		14'h15ad: data = 9'o152;
		14'h15ae: data = 9'o52;
		14'h15af: data = 9'o52;
		14'h15b0: data = 9'o152;
		14'h15b1: data = 9'o153;
		14'h15b2: data = 9'o52;
		14'h15b3: data = 9'o52;
		14'h15b4: data = 9'o162;
		14'h15b5: data = 9'o272;
		14'h15b6: data = 9'o172;
		14'h15b7: data = 9'o272;
		14'h15b8: data = 9'o372;
		14'h15b9: data = 9'o373;
		14'h15ba: data = 9'o273;
		14'h15bb: data = 9'o272;
		14'h15bc: data = 9'o272;
		14'h15bd: data = 9'o172;
		14'h15be: data = 9'o272;
		14'h15bf: data = 9'o272;
		14'h15c0: data = 9'o272;
		14'h15c1: data = 9'o172;
		14'h15c2: data = 9'o272;
		14'h15c3: data = 9'o272;
		14'h15c4: data = 9'o272;
		14'h15c5: data = 9'o272;
		14'h15c6: data = 9'o272;
		14'h15c7: data = 9'o273;
		14'h15c8: data = 9'o273;
		14'h15c9: data = 9'o272;
		14'h15ca: data = 9'o272;
		14'h15cb: data = 9'o272;
		14'h15cc: data = 9'o272;
		14'h15cd: data = 9'o272;
		14'h15ce: data = 9'o172;
		14'h15cf: data = 9'o172;
		14'h15d0: data = 9'o272;
		14'h15d1: data = 9'o473;
		14'h15d2: data = 9'o773;
		14'h15d3: data = 9'o773;
		14'h15d4: data = 9'o773;
		14'h15d5: data = 9'o762;
		14'h15d6: data = 9'o0;
		14'h15d7: data = 9'o0;
		14'h15d8: data = 9'o0;
		14'h15d9: data = 9'o0;
		14'h15da: data = 9'o0;
		14'h15db: data = 9'o0;
		14'h15dc: data = 9'o0;
		14'h15dd: data = 9'o0;
		14'h15de: data = 9'o0;
		14'h15df: data = 9'o0;
		14'h15e0: data = 9'o0;
		14'h15e1: data = 9'o0;
		14'h15e2: data = 9'o0;
		14'h15e3: data = 9'o0;
		14'h15e4: data = 9'o0;
		14'h15e5: data = 9'o0;
		14'h15e6: data = 9'o0;
		14'h15e7: data = 9'o651;
		14'h15e8: data = 9'o762;
		14'h15e9: data = 9'o773;
		14'h15ea: data = 9'o773;
		14'h15eb: data = 9'o673;
		14'h15ec: data = 9'o473;
		14'h15ed: data = 9'o272;
		14'h15ee: data = 9'o272;
		14'h15ef: data = 9'o172;
		14'h15f0: data = 9'o172;
		14'h15f1: data = 9'o172;
		14'h15f2: data = 9'o273;
		14'h15f3: data = 9'o272;
		14'h15f4: data = 9'o272;
		14'h15f5: data = 9'o172;
		14'h15f6: data = 9'o172;
		14'h15f7: data = 9'o272;
		14'h15f8: data = 9'o172;
		14'h15f9: data = 9'o172;
		14'h15fa: data = 9'o273;
		14'h15fb: data = 9'o172;
		14'h15fc: data = 9'o172;
		14'h15fd: data = 9'o172;
		14'h15fe: data = 9'o172;
		14'h15ff: data = 9'o172;
		14'h1600: data = 9'o272;
		14'h1601: data = 9'o272;
		14'h1602: data = 9'o272;
		14'h1603: data = 9'o172;
		14'h1604: data = 9'o273;
		14'h1605: data = 9'o272;
		14'h1606: data = 9'o272;
		14'h1607: data = 9'o272;
		14'h1608: data = 9'o273;
		14'h1609: data = 9'o172;
		14'h160a: data = 9'o52;
		14'h160b: data = 9'o152;
		14'h160c: data = 9'o52;
		14'h160d: data = 9'o152;
		14'h160e: data = 9'o52;
		14'h160f: data = 9'o52;
		14'h1610: data = 9'o52;
		14'h1611: data = 9'o152;
		14'h1612: data = 9'o52;
		14'h1613: data = 9'o52;
		14'h1614: data = 9'o152;
		14'h1615: data = 9'o152;
		14'h1616: data = 9'o52;
		14'h1617: data = 9'o52;
		14'h1618: data = 9'o162;
		14'h1619: data = 9'o272;
		14'h161a: data = 9'o172;
		14'h161b: data = 9'o172;
		14'h161c: data = 9'o272;
		14'h161d: data = 9'o272;
		14'h161e: data = 9'o273;
		14'h161f: data = 9'o172;
		14'h1620: data = 9'o272;
		14'h1621: data = 9'o172;
		14'h1622: data = 9'o272;
		14'h1623: data = 9'o172;
		14'h1624: data = 9'o172;
		14'h1625: data = 9'o172;
		14'h1626: data = 9'o172;
		14'h1627: data = 9'o172;
		14'h1628: data = 9'o172;
		14'h1629: data = 9'o172;
		14'h162a: data = 9'o172;
		14'h162b: data = 9'o172;
		14'h162c: data = 9'o273;
		14'h162d: data = 9'o172;
		14'h162e: data = 9'o172;
		14'h162f: data = 9'o272;
		14'h1630: data = 9'o272;
		14'h1631: data = 9'o172;
		14'h1632: data = 9'o172;
		14'h1633: data = 9'o172;
		14'h1634: data = 9'o272;
		14'h1635: data = 9'o373;
		14'h1636: data = 9'o773;
		14'h1637: data = 9'o773;
		14'h1638: data = 9'o773;
		14'h1639: data = 9'o762;
		14'h163a: data = 9'o0;
		14'h163b: data = 9'o0;
		14'h163c: data = 9'o0;
		14'h163d: data = 9'o0;
		14'h163e: data = 9'o0;
		14'h163f: data = 9'o0;
		14'h1640: data = 9'o0;
		14'h1641: data = 9'o0;
		14'h1642: data = 9'o0;
		14'h1643: data = 9'o0;
		14'h1644: data = 9'o0;
		14'h1645: data = 9'o0;
		14'h1646: data = 9'o0;
		14'h1647: data = 9'o0;
		14'h1648: data = 9'o0;
		14'h1649: data = 9'o0;
		14'h164a: data = 9'o0;
		14'h164b: data = 9'o651;
		14'h164c: data = 9'o762;
		14'h164d: data = 9'o773;
		14'h164e: data = 9'o773;
		14'h164f: data = 9'o773;
		14'h1650: data = 9'o372;
		14'h1651: data = 9'o272;
		14'h1652: data = 9'o172;
		14'h1653: data = 9'o172;
		14'h1654: data = 9'o172;
		14'h1655: data = 9'o172;
		14'h1656: data = 9'o272;
		14'h1657: data = 9'o272;
		14'h1658: data = 9'o172;
		14'h1659: data = 9'o172;
		14'h165a: data = 9'o172;
		14'h165b: data = 9'o172;
		14'h165c: data = 9'o172;
		14'h165d: data = 9'o172;
		14'h165e: data = 9'o172;
		14'h165f: data = 9'o172;
		14'h1660: data = 9'o172;
		14'h1661: data = 9'o172;
		14'h1662: data = 9'o172;
		14'h1663: data = 9'o172;
		14'h1664: data = 9'o172;
		14'h1665: data = 9'o172;
		14'h1666: data = 9'o272;
		14'h1667: data = 9'o172;
		14'h1668: data = 9'o273;
		14'h1669: data = 9'o273;
		14'h166a: data = 9'o272;
		14'h166b: data = 9'o272;
		14'h166c: data = 9'o273;
		14'h166d: data = 9'o162;
		14'h166e: data = 9'o152;
		14'h166f: data = 9'o152;
		14'h1670: data = 9'o152;
		14'h1671: data = 9'o52;
		14'h1672: data = 9'o52;
		14'h1673: data = 9'o52;
		14'h1674: data = 9'o52;
		14'h1675: data = 9'o52;
		14'h1676: data = 9'o52;
		14'h1677: data = 9'o152;
		14'h1678: data = 9'o152;
		14'h1679: data = 9'o152;
		14'h167a: data = 9'o52;
		14'h167b: data = 9'o52;
		14'h167c: data = 9'o162;
		14'h167d: data = 9'o273;
		14'h167e: data = 9'o172;
		14'h167f: data = 9'o172;
		14'h1680: data = 9'o273;
		14'h1681: data = 9'o272;
		14'h1682: data = 9'o273;
		14'h1683: data = 9'o273;
		14'h1684: data = 9'o172;
		14'h1685: data = 9'o172;
		14'h1686: data = 9'o172;
		14'h1687: data = 9'o172;
		14'h1688: data = 9'o172;
		14'h1689: data = 9'o172;
		14'h168a: data = 9'o172;
		14'h168b: data = 9'o172;
		14'h168c: data = 9'o172;
		14'h168d: data = 9'o172;
		14'h168e: data = 9'o172;
		14'h168f: data = 9'o172;
		14'h1690: data = 9'o172;
		14'h1691: data = 9'o172;
		14'h1692: data = 9'o172;
		14'h1693: data = 9'o172;
		14'h1694: data = 9'o172;
		14'h1695: data = 9'o172;
		14'h1696: data = 9'o172;
		14'h1697: data = 9'o172;
		14'h1698: data = 9'o172;
		14'h1699: data = 9'o372;
		14'h169a: data = 9'o773;
		14'h169b: data = 9'o773;
		14'h169c: data = 9'o773;
		14'h169d: data = 9'o662;
		14'h169e: data = 9'o0;
		14'h169f: data = 9'o0;
		14'h16a0: data = 9'o0;
		14'h16a1: data = 9'o0;
		14'h16a2: data = 9'o0;
		14'h16a3: data = 9'o0;
		14'h16a4: data = 9'o0;
		14'h16a5: data = 9'o0;
		14'h16a6: data = 9'o0;
		14'h16a7: data = 9'o0;
		14'h16a8: data = 9'o0;
		14'h16a9: data = 9'o0;
		14'h16aa: data = 9'o0;
		14'h16ab: data = 9'o0;
		14'h16ac: data = 9'o0;
		14'h16ad: data = 9'o0;
		14'h16ae: data = 9'o0;
		14'h16af: data = 9'o651;
		14'h16b0: data = 9'o763;
		14'h16b1: data = 9'o773;
		14'h16b2: data = 9'o773;
		14'h16b3: data = 9'o673;
		14'h16b4: data = 9'o272;
		14'h16b5: data = 9'o172;
		14'h16b6: data = 9'o172;
		14'h16b7: data = 9'o172;
		14'h16b8: data = 9'o172;
		14'h16b9: data = 9'o172;
		14'h16ba: data = 9'o172;
		14'h16bb: data = 9'o172;
		14'h16bc: data = 9'o172;
		14'h16bd: data = 9'o172;
		14'h16be: data = 9'o172;
		14'h16bf: data = 9'o172;
		14'h16c0: data = 9'o172;
		14'h16c1: data = 9'o172;
		14'h16c2: data = 9'o172;
		14'h16c3: data = 9'o172;
		14'h16c4: data = 9'o172;
		14'h16c5: data = 9'o172;
		14'h16c6: data = 9'o172;
		14'h16c7: data = 9'o172;
		14'h16c8: data = 9'o172;
		14'h16c9: data = 9'o172;
		14'h16ca: data = 9'o273;
		14'h16cb: data = 9'o172;
		14'h16cc: data = 9'o273;
		14'h16cd: data = 9'o273;
		14'h16ce: data = 9'o172;
		14'h16cf: data = 9'o172;
		14'h16d0: data = 9'o272;
		14'h16d1: data = 9'o162;
		14'h16d2: data = 9'o152;
		14'h16d3: data = 9'o152;
		14'h16d4: data = 9'o152;
		14'h16d5: data = 9'o152;
		14'h16d6: data = 9'o52;
		14'h16d7: data = 9'o52;
		14'h16d8: data = 9'o52;
		14'h16d9: data = 9'o52;
		14'h16da: data = 9'o52;
		14'h16db: data = 9'o152;
		14'h16dc: data = 9'o152;
		14'h16dd: data = 9'o152;
		14'h16de: data = 9'o152;
		14'h16df: data = 9'o52;
		14'h16e0: data = 9'o162;
		14'h16e1: data = 9'o173;
		14'h16e2: data = 9'o172;
		14'h16e3: data = 9'o172;
		14'h16e4: data = 9'o273;
		14'h16e5: data = 9'o273;
		14'h16e6: data = 9'o172;
		14'h16e7: data = 9'o272;
		14'h16e8: data = 9'o172;
		14'h16e9: data = 9'o172;
		14'h16ea: data = 9'o172;
		14'h16eb: data = 9'o172;
		14'h16ec: data = 9'o172;
		14'h16ed: data = 9'o172;
		14'h16ee: data = 9'o172;
		14'h16ef: data = 9'o172;
		14'h16f0: data = 9'o172;
		14'h16f1: data = 9'o172;
		14'h16f2: data = 9'o172;
		14'h16f3: data = 9'o172;
		14'h16f4: data = 9'o172;
		14'h16f5: data = 9'o172;
		14'h16f6: data = 9'o172;
		14'h16f7: data = 9'o172;
		14'h16f8: data = 9'o172;
		14'h16f9: data = 9'o172;
		14'h16fa: data = 9'o172;
		14'h16fb: data = 9'o172;
		14'h16fc: data = 9'o172;
		14'h16fd: data = 9'o272;
		14'h16fe: data = 9'o673;
		14'h16ff: data = 9'o773;
		14'h1700: data = 9'o773;
		14'h1701: data = 9'o662;
		14'h1702: data = 9'o0;
		14'h1703: data = 9'o0;
		14'h1704: data = 9'o0;
		14'h1705: data = 9'o0;
		14'h1706: data = 9'o0;
		14'h1707: data = 9'o0;
		14'h1708: data = 9'o0;
		14'h1709: data = 9'o0;
		14'h170a: data = 9'o0;
		14'h170b: data = 9'o0;
		14'h170c: data = 9'o0;
		14'h170d: data = 9'o0;
		14'h170e: data = 9'o0;
		14'h170f: data = 9'o0;
		14'h1710: data = 9'o0;
		14'h1711: data = 9'o0;
		14'h1712: data = 9'o0;
		14'h1713: data = 9'o651;
		14'h1714: data = 9'o762;
		14'h1715: data = 9'o773;
		14'h1716: data = 9'o773;
		14'h1717: data = 9'o673;
		14'h1718: data = 9'o272;
		14'h1719: data = 9'o172;
		14'h171a: data = 9'o172;
		14'h171b: data = 9'o172;
		14'h171c: data = 9'o172;
		14'h171d: data = 9'o172;
		14'h171e: data = 9'o172;
		14'h171f: data = 9'o172;
		14'h1720: data = 9'o172;
		14'h1721: data = 9'o172;
		14'h1722: data = 9'o172;
		14'h1723: data = 9'o172;
		14'h1724: data = 9'o172;
		14'h1725: data = 9'o172;
		14'h1726: data = 9'o172;
		14'h1727: data = 9'o172;
		14'h1728: data = 9'o172;
		14'h1729: data = 9'o172;
		14'h172a: data = 9'o172;
		14'h172b: data = 9'o172;
		14'h172c: data = 9'o172;
		14'h172d: data = 9'o172;
		14'h172e: data = 9'o272;
		14'h172f: data = 9'o162;
		14'h1730: data = 9'o162;
		14'h1731: data = 9'o162;
		14'h1732: data = 9'o172;
		14'h1733: data = 9'o272;
		14'h1734: data = 9'o273;
		14'h1735: data = 9'o172;
		14'h1736: data = 9'o52;
		14'h1737: data = 9'o52;
		14'h1738: data = 9'o152;
		14'h1739: data = 9'o152;
		14'h173a: data = 9'o52;
		14'h173b: data = 9'o52;
		14'h173c: data = 9'o52;
		14'h173d: data = 9'o52;
		14'h173e: data = 9'o152;
		14'h173f: data = 9'o152;
		14'h1740: data = 9'o152;
		14'h1741: data = 9'o152;
		14'h1742: data = 9'o52;
		14'h1743: data = 9'o52;
		14'h1744: data = 9'o162;
		14'h1745: data = 9'o273;
		14'h1746: data = 9'o273;
		14'h1747: data = 9'o173;
		14'h1748: data = 9'o162;
		14'h1749: data = 9'o62;
		14'h174a: data = 9'o162;
		14'h174b: data = 9'o172;
		14'h174c: data = 9'o172;
		14'h174d: data = 9'o172;
		14'h174e: data = 9'o172;
		14'h174f: data = 9'o172;
		14'h1750: data = 9'o172;
		14'h1751: data = 9'o172;
		14'h1752: data = 9'o172;
		14'h1753: data = 9'o172;
		14'h1754: data = 9'o172;
		14'h1755: data = 9'o172;
		14'h1756: data = 9'o172;
		14'h1757: data = 9'o172;
		14'h1758: data = 9'o172;
		14'h1759: data = 9'o172;
		14'h175a: data = 9'o172;
		14'h175b: data = 9'o172;
		14'h175c: data = 9'o172;
		14'h175d: data = 9'o172;
		14'h175e: data = 9'o172;
		14'h175f: data = 9'o172;
		14'h1760: data = 9'o172;
		14'h1761: data = 9'o272;
		14'h1762: data = 9'o673;
		14'h1763: data = 9'o773;
		14'h1764: data = 9'o773;
		14'h1765: data = 9'o662;
		14'h1766: data = 9'o0;
		14'h1767: data = 9'o0;
		14'h1768: data = 9'o0;
		14'h1769: data = 9'o0;
		14'h176a: data = 9'o0;
		14'h176b: data = 9'o0;
		14'h176c: data = 9'o0;
		14'h176d: data = 9'o0;
		14'h176e: data = 9'o0;
		14'h176f: data = 9'o0;
		14'h1770: data = 9'o0;
		14'h1771: data = 9'o0;
		14'h1772: data = 9'o0;
		14'h1773: data = 9'o0;
		14'h1774: data = 9'o0;
		14'h1775: data = 9'o0;
		14'h1776: data = 9'o0;
		14'h1777: data = 9'o651;
		14'h1778: data = 9'o762;
		14'h1779: data = 9'o773;
		14'h177a: data = 9'o773;
		14'h177b: data = 9'o673;
		14'h177c: data = 9'o272;
		14'h177d: data = 9'o172;
		14'h177e: data = 9'o172;
		14'h177f: data = 9'o172;
		14'h1780: data = 9'o172;
		14'h1781: data = 9'o172;
		14'h1782: data = 9'o172;
		14'h1783: data = 9'o172;
		14'h1784: data = 9'o172;
		14'h1785: data = 9'o172;
		14'h1786: data = 9'o172;
		14'h1787: data = 9'o172;
		14'h1788: data = 9'o172;
		14'h1789: data = 9'o172;
		14'h178a: data = 9'o172;
		14'h178b: data = 9'o172;
		14'h178c: data = 9'o172;
		14'h178d: data = 9'o172;
		14'h178e: data = 9'o172;
		14'h178f: data = 9'o172;
		14'h1790: data = 9'o172;
		14'h1791: data = 9'o172;
		14'h1792: data = 9'o172;
		14'h1793: data = 9'o62;
		14'h1794: data = 9'o52;
		14'h1795: data = 9'o52;
		14'h1796: data = 9'o172;
		14'h1797: data = 9'o172;
		14'h1798: data = 9'o173;
		14'h1799: data = 9'o172;
		14'h179a: data = 9'o52;
		14'h179b: data = 9'o52;
		14'h179c: data = 9'o152;
		14'h179d: data = 9'o152;
		14'h179e: data = 9'o152;
		14'h179f: data = 9'o152;
		14'h17a0: data = 9'o52;
		14'h17a1: data = 9'o152;
		14'h17a2: data = 9'o152;
		14'h17a3: data = 9'o152;
		14'h17a4: data = 9'o152;
		14'h17a5: data = 9'o152;
		14'h17a6: data = 9'o152;
		14'h17a7: data = 9'o52;
		14'h17a8: data = 9'o173;
		14'h17a9: data = 9'o273;
		14'h17aa: data = 9'o273;
		14'h17ab: data = 9'o273;
		14'h17ac: data = 9'o62;
		14'h17ad: data = 9'o52;
		14'h17ae: data = 9'o52;
		14'h17af: data = 9'o172;
		14'h17b0: data = 9'o272;
		14'h17b1: data = 9'o172;
		14'h17b2: data = 9'o172;
		14'h17b3: data = 9'o172;
		14'h17b4: data = 9'o272;
		14'h17b5: data = 9'o172;
		14'h17b6: data = 9'o172;
		14'h17b7: data = 9'o172;
		14'h17b8: data = 9'o172;
		14'h17b9: data = 9'o172;
		14'h17ba: data = 9'o172;
		14'h17bb: data = 9'o172;
		14'h17bc: data = 9'o172;
		14'h17bd: data = 9'o172;
		14'h17be: data = 9'o172;
		14'h17bf: data = 9'o172;
		14'h17c0: data = 9'o172;
		14'h17c1: data = 9'o172;
		14'h17c2: data = 9'o172;
		14'h17c3: data = 9'o172;
		14'h17c4: data = 9'o172;
		14'h17c5: data = 9'o272;
		14'h17c6: data = 9'o673;
		14'h17c7: data = 9'o773;
		14'h17c8: data = 9'o773;
		14'h17c9: data = 9'o763;
		14'h17ca: data = 9'o0;
		14'h17cb: data = 9'o0;
		14'h17cc: data = 9'o0;
		14'h17cd: data = 9'o0;
		14'h17ce: data = 9'o0;
		14'h17cf: data = 9'o0;
		14'h17d0: data = 9'o0;
		14'h17d1: data = 9'o0;
		14'h17d2: data = 9'o0;
		14'h17d3: data = 9'o0;
		14'h17d4: data = 9'o0;
		14'h17d5: data = 9'o0;
		14'h17d6: data = 9'o0;
		14'h17d7: data = 9'o0;
		14'h17d8: data = 9'o0;
		14'h17d9: data = 9'o0;
		14'h17da: data = 9'o0;
		14'h17db: data = 9'o651;
		14'h17dc: data = 9'o762;
		14'h17dd: data = 9'o773;
		14'h17de: data = 9'o773;
		14'h17df: data = 9'o573;
		14'h17e0: data = 9'o272;
		14'h17e1: data = 9'o172;
		14'h17e2: data = 9'o172;
		14'h17e3: data = 9'o172;
		14'h17e4: data = 9'o172;
		14'h17e5: data = 9'o172;
		14'h17e6: data = 9'o172;
		14'h17e7: data = 9'o172;
		14'h17e8: data = 9'o172;
		14'h17e9: data = 9'o172;
		14'h17ea: data = 9'o172;
		14'h17eb: data = 9'o172;
		14'h17ec: data = 9'o172;
		14'h17ed: data = 9'o172;
		14'h17ee: data = 9'o172;
		14'h17ef: data = 9'o172;
		14'h17f0: data = 9'o172;
		14'h17f1: data = 9'o172;
		14'h17f2: data = 9'o172;
		14'h17f3: data = 9'o172;
		14'h17f4: data = 9'o172;
		14'h17f5: data = 9'o272;
		14'h17f6: data = 9'o172;
		14'h17f7: data = 9'o52;
		14'h17f8: data = 9'o52;
		14'h17f9: data = 9'o62;
		14'h17fa: data = 9'o273;
		14'h17fb: data = 9'o273;
		14'h17fc: data = 9'o273;
		14'h17fd: data = 9'o173;
		14'h17fe: data = 9'o52;
		14'h17ff: data = 9'o52;
		14'h1800: data = 9'o52;
		14'h1801: data = 9'o152;
		14'h1802: data = 9'o152;
		14'h1803: data = 9'o152;
		14'h1804: data = 9'o152;
		14'h1805: data = 9'o152;
		14'h1806: data = 9'o152;
		14'h1807: data = 9'o152;
		14'h1808: data = 9'o152;
		14'h1809: data = 9'o52;
		14'h180a: data = 9'o152;
		14'h180b: data = 9'o52;
		14'h180c: data = 9'o163;
		14'h180d: data = 9'o273;
		14'h180e: data = 9'o273;
		14'h180f: data = 9'o273;
		14'h1810: data = 9'o52;
		14'h1811: data = 9'o52;
		14'h1812: data = 9'o52;
		14'h1813: data = 9'o272;
		14'h1814: data = 9'o273;
		14'h1815: data = 9'o172;
		14'h1816: data = 9'o172;
		14'h1817: data = 9'o172;
		14'h1818: data = 9'o172;
		14'h1819: data = 9'o172;
		14'h181a: data = 9'o172;
		14'h181b: data = 9'o172;
		14'h181c: data = 9'o172;
		14'h181d: data = 9'o172;
		14'h181e: data = 9'o172;
		14'h181f: data = 9'o172;
		14'h1820: data = 9'o172;
		14'h1821: data = 9'o172;
		14'h1822: data = 9'o172;
		14'h1823: data = 9'o172;
		14'h1824: data = 9'o172;
		14'h1825: data = 9'o172;
		14'h1826: data = 9'o172;
		14'h1827: data = 9'o172;
		14'h1828: data = 9'o172;
		14'h1829: data = 9'o272;
		14'h182a: data = 9'o573;
		14'h182b: data = 9'o773;
		14'h182c: data = 9'o773;
		14'h182d: data = 9'o763;
		14'h182e: data = 9'o0;
		14'h182f: data = 9'o0;
		14'h1830: data = 9'o0;
		14'h1831: data = 9'o0;
		14'h1832: data = 9'o0;
		14'h1833: data = 9'o0;
		14'h1834: data = 9'o0;
		14'h1835: data = 9'o0;
		14'h1836: data = 9'o0;
		14'h1837: data = 9'o0;
		14'h1838: data = 9'o0;
		14'h1839: data = 9'o0;
		14'h183a: data = 9'o0;
		14'h183b: data = 9'o0;
		14'h183c: data = 9'o0;
		14'h183d: data = 9'o0;
		14'h183e: data = 9'o0;
		14'h183f: data = 9'o651;
		14'h1840: data = 9'o762;
		14'h1841: data = 9'o773;
		14'h1842: data = 9'o773;
		14'h1843: data = 9'o573;
		14'h1844: data = 9'o272;
		14'h1845: data = 9'o172;
		14'h1846: data = 9'o272;
		14'h1847: data = 9'o172;
		14'h1848: data = 9'o172;
		14'h1849: data = 9'o172;
		14'h184a: data = 9'o172;
		14'h184b: data = 9'o172;
		14'h184c: data = 9'o172;
		14'h184d: data = 9'o172;
		14'h184e: data = 9'o172;
		14'h184f: data = 9'o172;
		14'h1850: data = 9'o172;
		14'h1851: data = 9'o172;
		14'h1852: data = 9'o172;
		14'h1853: data = 9'o172;
		14'h1854: data = 9'o172;
		14'h1855: data = 9'o172;
		14'h1856: data = 9'o172;
		14'h1857: data = 9'o172;
		14'h1858: data = 9'o172;
		14'h1859: data = 9'o272;
		14'h185a: data = 9'o273;
		14'h185b: data = 9'o52;
		14'h185c: data = 9'o52;
		14'h185d: data = 9'o52;
		14'h185e: data = 9'o273;
		14'h185f: data = 9'o273;
		14'h1860: data = 9'o273;
		14'h1861: data = 9'o163;
		14'h1862: data = 9'o52;
		14'h1863: data = 9'o52;
		14'h1864: data = 9'o52;
		14'h1865: data = 9'o152;
		14'h1866: data = 9'o152;
		14'h1867: data = 9'o152;
		14'h1868: data = 9'o152;
		14'h1869: data = 9'o152;
		14'h186a: data = 9'o152;
		14'h186b: data = 9'o52;
		14'h186c: data = 9'o52;
		14'h186d: data = 9'o52;
		14'h186e: data = 9'o152;
		14'h186f: data = 9'o152;
		14'h1870: data = 9'o163;
		14'h1871: data = 9'o273;
		14'h1872: data = 9'o273;
		14'h1873: data = 9'o273;
		14'h1874: data = 9'o162;
		14'h1875: data = 9'o52;
		14'h1876: data = 9'o52;
		14'h1877: data = 9'o273;
		14'h1878: data = 9'o273;
		14'h1879: data = 9'o172;
		14'h187a: data = 9'o172;
		14'h187b: data = 9'o172;
		14'h187c: data = 9'o172;
		14'h187d: data = 9'o172;
		14'h187e: data = 9'o172;
		14'h187f: data = 9'o172;
		14'h1880: data = 9'o172;
		14'h1881: data = 9'o172;
		14'h1882: data = 9'o172;
		14'h1883: data = 9'o172;
		14'h1884: data = 9'o172;
		14'h1885: data = 9'o172;
		14'h1886: data = 9'o172;
		14'h1887: data = 9'o172;
		14'h1888: data = 9'o172;
		14'h1889: data = 9'o172;
		14'h188a: data = 9'o172;
		14'h188b: data = 9'o172;
		14'h188c: data = 9'o172;
		14'h188d: data = 9'o272;
		14'h188e: data = 9'o573;
		14'h188f: data = 9'o773;
		14'h1890: data = 9'o773;
		14'h1891: data = 9'o662;
		14'h1892: data = 9'o0;
		14'h1893: data = 9'o0;
		14'h1894: data = 9'o0;
		14'h1895: data = 9'o0;
		14'h1896: data = 9'o0;
		14'h1897: data = 9'o0;
		14'h1898: data = 9'o0;
		14'h1899: data = 9'o0;
		14'h189a: data = 9'o0;
		14'h189b: data = 9'o0;
		14'h189c: data = 9'o0;
		14'h189d: data = 9'o0;
		14'h189e: data = 9'o0;
		14'h189f: data = 9'o0;
		14'h18a0: data = 9'o0;
		14'h18a1: data = 9'o0;
		14'h18a2: data = 9'o0;
		14'h18a3: data = 9'o651;
		14'h18a4: data = 9'o762;
		14'h18a5: data = 9'o773;
		14'h18a6: data = 9'o773;
		14'h18a7: data = 9'o473;
		14'h18a8: data = 9'o272;
		14'h18a9: data = 9'o172;
		14'h18aa: data = 9'o272;
		14'h18ab: data = 9'o172;
		14'h18ac: data = 9'o172;
		14'h18ad: data = 9'o172;
		14'h18ae: data = 9'o172;
		14'h18af: data = 9'o172;
		14'h18b0: data = 9'o172;
		14'h18b1: data = 9'o172;
		14'h18b2: data = 9'o172;
		14'h18b3: data = 9'o172;
		14'h18b4: data = 9'o172;
		14'h18b5: data = 9'o172;
		14'h18b6: data = 9'o172;
		14'h18b7: data = 9'o172;
		14'h18b8: data = 9'o172;
		14'h18b9: data = 9'o172;
		14'h18ba: data = 9'o172;
		14'h18bb: data = 9'o172;
		14'h18bc: data = 9'o272;
		14'h18bd: data = 9'o272;
		14'h18be: data = 9'o273;
		14'h18bf: data = 9'o52;
		14'h18c0: data = 9'o52;
		14'h18c1: data = 9'o52;
		14'h18c2: data = 9'o52;
		14'h18c3: data = 9'o52;
		14'h18c4: data = 9'o52;
		14'h18c5: data = 9'o152;
		14'h18c6: data = 9'o52;
		14'h18c7: data = 9'o52;
		14'h18c8: data = 9'o152;
		14'h18c9: data = 9'o152;
		14'h18ca: data = 9'o152;
		14'h18cb: data = 9'o152;
		14'h18cc: data = 9'o152;
		14'h18cd: data = 9'o152;
		14'h18ce: data = 9'o152;
		14'h18cf: data = 9'o52;
		14'h18d0: data = 9'o52;
		14'h18d1: data = 9'o52;
		14'h18d2: data = 9'o152;
		14'h18d3: data = 9'o52;
		14'h18d4: data = 9'o52;
		14'h18d5: data = 9'o52;
		14'h18d6: data = 9'o52;
		14'h18d7: data = 9'o52;
		14'h18d8: data = 9'o52;
		14'h18d9: data = 9'o52;
		14'h18da: data = 9'o52;
		14'h18db: data = 9'o273;
		14'h18dc: data = 9'o272;
		14'h18dd: data = 9'o172;
		14'h18de: data = 9'o172;
		14'h18df: data = 9'o172;
		14'h18e0: data = 9'o172;
		14'h18e1: data = 9'o272;
		14'h18e2: data = 9'o172;
		14'h18e3: data = 9'o172;
		14'h18e4: data = 9'o172;
		14'h18e5: data = 9'o172;
		14'h18e6: data = 9'o172;
		14'h18e7: data = 9'o172;
		14'h18e8: data = 9'o172;
		14'h18e9: data = 9'o172;
		14'h18ea: data = 9'o172;
		14'h18eb: data = 9'o172;
		14'h18ec: data = 9'o172;
		14'h18ed: data = 9'o172;
		14'h18ee: data = 9'o172;
		14'h18ef: data = 9'o172;
		14'h18f0: data = 9'o172;
		14'h18f1: data = 9'o272;
		14'h18f2: data = 9'o473;
		14'h18f3: data = 9'o773;
		14'h18f4: data = 9'o773;
		14'h18f5: data = 9'o762;
		14'h18f6: data = 9'o0;
		14'h18f7: data = 9'o0;
		14'h18f8: data = 9'o0;
		14'h18f9: data = 9'o0;
		14'h18fa: data = 9'o0;
		14'h18fb: data = 9'o0;
		14'h18fc: data = 9'o0;
		14'h18fd: data = 9'o0;
		14'h18fe: data = 9'o0;
		14'h18ff: data = 9'o0;
		14'h1900: data = 9'o0;
		14'h1901: data = 9'o0;
		14'h1902: data = 9'o0;
		14'h1903: data = 9'o0;
		14'h1904: data = 9'o0;
		14'h1905: data = 9'o0;
		14'h1906: data = 9'o0;
		14'h1907: data = 9'o652;
		14'h1908: data = 9'o762;
		14'h1909: data = 9'o773;
		14'h190a: data = 9'o673;
		14'h190b: data = 9'o473;
		14'h190c: data = 9'o272;
		14'h190d: data = 9'o172;
		14'h190e: data = 9'o272;
		14'h190f: data = 9'o172;
		14'h1910: data = 9'o172;
		14'h1911: data = 9'o172;
		14'h1912: data = 9'o172;
		14'h1913: data = 9'o172;
		14'h1914: data = 9'o172;
		14'h1915: data = 9'o172;
		14'h1916: data = 9'o172;
		14'h1917: data = 9'o172;
		14'h1918: data = 9'o172;
		14'h1919: data = 9'o172;
		14'h191a: data = 9'o172;
		14'h191b: data = 9'o172;
		14'h191c: data = 9'o172;
		14'h191d: data = 9'o172;
		14'h191e: data = 9'o172;
		14'h191f: data = 9'o172;
		14'h1920: data = 9'o272;
		14'h1921: data = 9'o273;
		14'h1922: data = 9'o273;
		14'h1923: data = 9'o52;
		14'h1924: data = 9'o52;
		14'h1925: data = 9'o152;
		14'h1926: data = 9'o152;
		14'h1927: data = 9'o52;
		14'h1928: data = 9'o52;
		14'h1929: data = 9'o152;
		14'h192a: data = 9'o52;
		14'h192b: data = 9'o152;
		14'h192c: data = 9'o152;
		14'h192d: data = 9'o152;
		14'h192e: data = 9'o152;
		14'h192f: data = 9'o152;
		14'h1930: data = 9'o152;
		14'h1931: data = 9'o152;
		14'h1932: data = 9'o152;
		14'h1933: data = 9'o152;
		14'h1934: data = 9'o52;
		14'h1935: data = 9'o52;
		14'h1936: data = 9'o152;
		14'h1937: data = 9'o152;
		14'h1938: data = 9'o52;
		14'h1939: data = 9'o52;
		14'h193a: data = 9'o52;
		14'h193b: data = 9'o52;
		14'h193c: data = 9'o52;
		14'h193d: data = 9'o52;
		14'h193e: data = 9'o52;
		14'h193f: data = 9'o273;
		14'h1940: data = 9'o272;
		14'h1941: data = 9'o172;
		14'h1942: data = 9'o272;
		14'h1943: data = 9'o172;
		14'h1944: data = 9'o172;
		14'h1945: data = 9'o172;
		14'h1946: data = 9'o172;
		14'h1947: data = 9'o172;
		14'h1948: data = 9'o172;
		14'h1949: data = 9'o172;
		14'h194a: data = 9'o172;
		14'h194b: data = 9'o172;
		14'h194c: data = 9'o172;
		14'h194d: data = 9'o172;
		14'h194e: data = 9'o172;
		14'h194f: data = 9'o172;
		14'h1950: data = 9'o172;
		14'h1951: data = 9'o172;
		14'h1952: data = 9'o172;
		14'h1953: data = 9'o172;
		14'h1954: data = 9'o172;
		14'h1955: data = 9'o272;
		14'h1956: data = 9'o473;
		14'h1957: data = 9'o673;
		14'h1958: data = 9'o773;
		14'h1959: data = 9'o763;
		14'h195a: data = 9'o0;
		14'h195b: data = 9'o0;
		14'h195c: data = 9'o0;
		14'h195d: data = 9'o0;
		14'h195e: data = 9'o0;
		14'h195f: data = 9'o0;
		14'h1960: data = 9'o0;
		14'h1961: data = 9'o0;
		14'h1962: data = 9'o0;
		14'h1963: data = 9'o0;
		14'h1964: data = 9'o0;
		14'h1965: data = 9'o0;
		14'h1966: data = 9'o0;
		14'h1967: data = 9'o0;
		14'h1968: data = 9'o0;
		14'h1969: data = 9'o0;
		14'h196a: data = 9'o0;
		14'h196b: data = 9'o651;
		14'h196c: data = 9'o662;
		14'h196d: data = 9'o773;
		14'h196e: data = 9'o673;
		14'h196f: data = 9'o373;
		14'h1970: data = 9'o272;
		14'h1971: data = 9'o172;
		14'h1972: data = 9'o272;
		14'h1973: data = 9'o172;
		14'h1974: data = 9'o172;
		14'h1975: data = 9'o172;
		14'h1976: data = 9'o172;
		14'h1977: data = 9'o172;
		14'h1978: data = 9'o172;
		14'h1979: data = 9'o172;
		14'h197a: data = 9'o172;
		14'h197b: data = 9'o172;
		14'h197c: data = 9'o172;
		14'h197d: data = 9'o172;
		14'h197e: data = 9'o172;
		14'h197f: data = 9'o172;
		14'h1980: data = 9'o172;
		14'h1981: data = 9'o172;
		14'h1982: data = 9'o172;
		14'h1983: data = 9'o172;
		14'h1984: data = 9'o172;
		14'h1985: data = 9'o273;
		14'h1986: data = 9'o273;
		14'h1987: data = 9'o52;
		14'h1988: data = 9'o52;
		14'h1989: data = 9'o152;
		14'h198a: data = 9'o52;
		14'h198b: data = 9'o152;
		14'h198c: data = 9'o152;
		14'h198d: data = 9'o52;
		14'h198e: data = 9'o152;
		14'h198f: data = 9'o152;
		14'h1990: data = 9'o152;
		14'h1991: data = 9'o252;
		14'h1992: data = 9'o142;
		14'h1993: data = 9'o142;
		14'h1994: data = 9'o142;
		14'h1995: data = 9'o142;
		14'h1996: data = 9'o152;
		14'h1997: data = 9'o152;
		14'h1998: data = 9'o152;
		14'h1999: data = 9'o152;
		14'h199a: data = 9'o152;
		14'h199b: data = 9'o142;
		14'h199c: data = 9'o152;
		14'h199d: data = 9'o152;
		14'h199e: data = 9'o52;
		14'h199f: data = 9'o52;
		14'h19a0: data = 9'o152;
		14'h19a1: data = 9'o52;
		14'h19a2: data = 9'o52;
		14'h19a3: data = 9'o273;
		14'h19a4: data = 9'o273;
		14'h19a5: data = 9'o172;
		14'h19a6: data = 9'o172;
		14'h19a7: data = 9'o172;
		14'h19a8: data = 9'o172;
		14'h19a9: data = 9'o172;
		14'h19aa: data = 9'o172;
		14'h19ab: data = 9'o172;
		14'h19ac: data = 9'o172;
		14'h19ad: data = 9'o172;
		14'h19ae: data = 9'o172;
		14'h19af: data = 9'o172;
		14'h19b0: data = 9'o172;
		14'h19b1: data = 9'o172;
		14'h19b2: data = 9'o172;
		14'h19b3: data = 9'o172;
		14'h19b4: data = 9'o172;
		14'h19b5: data = 9'o172;
		14'h19b6: data = 9'o172;
		14'h19b7: data = 9'o172;
		14'h19b8: data = 9'o172;
		14'h19b9: data = 9'o272;
		14'h19ba: data = 9'o372;
		14'h19bb: data = 9'o673;
		14'h19bc: data = 9'o773;
		14'h19bd: data = 9'o763;
		14'h19be: data = 9'o0;
		14'h19bf: data = 9'o0;
		14'h19c0: data = 9'o0;
		14'h19c1: data = 9'o0;
		14'h19c2: data = 9'o0;
		14'h19c3: data = 9'o0;
		14'h19c4: data = 9'o0;
		14'h19c5: data = 9'o0;
		14'h19c6: data = 9'o0;
		14'h19c7: data = 9'o0;
		14'h19c8: data = 9'o0;
		14'h19c9: data = 9'o0;
		14'h19ca: data = 9'o0;
		14'h19cb: data = 9'o0;
		14'h19cc: data = 9'o0;
		14'h19cd: data = 9'o0;
		14'h19ce: data = 9'o0;
		14'h19cf: data = 9'o651;
		14'h19d0: data = 9'o662;
		14'h19d1: data = 9'o773;
		14'h19d2: data = 9'o673;
		14'h19d3: data = 9'o373;
		14'h19d4: data = 9'o272;
		14'h19d5: data = 9'o172;
		14'h19d6: data = 9'o272;
		14'h19d7: data = 9'o172;
		14'h19d8: data = 9'o172;
		14'h19d9: data = 9'o172;
		14'h19da: data = 9'o172;
		14'h19db: data = 9'o172;
		14'h19dc: data = 9'o172;
		14'h19dd: data = 9'o172;
		14'h19de: data = 9'o172;
		14'h19df: data = 9'o172;
		14'h19e0: data = 9'o172;
		14'h19e1: data = 9'o172;
		14'h19e2: data = 9'o172;
		14'h19e3: data = 9'o172;
		14'h19e4: data = 9'o172;
		14'h19e5: data = 9'o172;
		14'h19e6: data = 9'o172;
		14'h19e7: data = 9'o172;
		14'h19e8: data = 9'o172;
		14'h19e9: data = 9'o273;
		14'h19ea: data = 9'o273;
		14'h19eb: data = 9'o52;
		14'h19ec: data = 9'o52;
		14'h19ed: data = 9'o152;
		14'h19ee: data = 9'o152;
		14'h19ef: data = 9'o152;
		14'h19f0: data = 9'o152;
		14'h19f1: data = 9'o152;
		14'h19f2: data = 9'o152;
		14'h19f3: data = 9'o152;
		14'h19f4: data = 9'o142;
		14'h19f5: data = 9'o31;
		14'h19f6: data = 9'o21;
		14'h19f7: data = 9'o21;
		14'h19f8: data = 9'o21;
		14'h19f9: data = 9'o21;
		14'h19fa: data = 9'o21;
		14'h19fb: data = 9'o31;
		14'h19fc: data = 9'o31;
		14'h19fd: data = 9'o142;
		14'h19fe: data = 9'o142;
		14'h19ff: data = 9'o152;
		14'h1a00: data = 9'o152;
		14'h1a01: data = 9'o52;
		14'h1a02: data = 9'o152;
		14'h1a03: data = 9'o52;
		14'h1a04: data = 9'o52;
		14'h1a05: data = 9'o52;
		14'h1a06: data = 9'o52;
		14'h1a07: data = 9'o273;
		14'h1a08: data = 9'o273;
		14'h1a09: data = 9'o172;
		14'h1a0a: data = 9'o172;
		14'h1a0b: data = 9'o172;
		14'h1a0c: data = 9'o172;
		14'h1a0d: data = 9'o172;
		14'h1a0e: data = 9'o172;
		14'h1a0f: data = 9'o172;
		14'h1a10: data = 9'o172;
		14'h1a11: data = 9'o172;
		14'h1a12: data = 9'o172;
		14'h1a13: data = 9'o172;
		14'h1a14: data = 9'o172;
		14'h1a15: data = 9'o172;
		14'h1a16: data = 9'o172;
		14'h1a17: data = 9'o172;
		14'h1a18: data = 9'o172;
		14'h1a19: data = 9'o172;
		14'h1a1a: data = 9'o172;
		14'h1a1b: data = 9'o172;
		14'h1a1c: data = 9'o172;
		14'h1a1d: data = 9'o272;
		14'h1a1e: data = 9'o372;
		14'h1a1f: data = 9'o673;
		14'h1a20: data = 9'o773;
		14'h1a21: data = 9'o762;
		14'h1a22: data = 9'o0;
		14'h1a23: data = 9'o0;
		14'h1a24: data = 9'o0;
		14'h1a25: data = 9'o0;
		14'h1a26: data = 9'o0;
		14'h1a27: data = 9'o0;
		14'h1a28: data = 9'o0;
		14'h1a29: data = 9'o0;
		14'h1a2a: data = 9'o0;
		14'h1a2b: data = 9'o0;
		14'h1a2c: data = 9'o0;
		14'h1a2d: data = 9'o0;
		14'h1a2e: data = 9'o0;
		14'h1a2f: data = 9'o0;
		14'h1a30: data = 9'o0;
		14'h1a31: data = 9'o0;
		14'h1a32: data = 9'o0;
		14'h1a33: data = 9'o651;
		14'h1a34: data = 9'o662;
		14'h1a35: data = 9'o773;
		14'h1a36: data = 9'o673;
		14'h1a37: data = 9'o372;
		14'h1a38: data = 9'o272;
		14'h1a39: data = 9'o172;
		14'h1a3a: data = 9'o172;
		14'h1a3b: data = 9'o172;
		14'h1a3c: data = 9'o172;
		14'h1a3d: data = 9'o172;
		14'h1a3e: data = 9'o172;
		14'h1a3f: data = 9'o172;
		14'h1a40: data = 9'o172;
		14'h1a41: data = 9'o172;
		14'h1a42: data = 9'o172;
		14'h1a43: data = 9'o172;
		14'h1a44: data = 9'o172;
		14'h1a45: data = 9'o172;
		14'h1a46: data = 9'o172;
		14'h1a47: data = 9'o172;
		14'h1a48: data = 9'o172;
		14'h1a49: data = 9'o172;
		14'h1a4a: data = 9'o172;
		14'h1a4b: data = 9'o172;
		14'h1a4c: data = 9'o172;
		14'h1a4d: data = 9'o273;
		14'h1a4e: data = 9'o273;
		14'h1a4f: data = 9'o52;
		14'h1a50: data = 9'o52;
		14'h1a51: data = 9'o52;
		14'h1a52: data = 9'o152;
		14'h1a53: data = 9'o52;
		14'h1a54: data = 9'o152;
		14'h1a55: data = 9'o152;
		14'h1a56: data = 9'o142;
		14'h1a57: data = 9'o32;
		14'h1a58: data = 9'o21;
		14'h1a59: data = 9'o21;
		14'h1a5a: data = 9'o11;
		14'h1a5b: data = 9'o10;
		14'h1a5c: data = 9'o10;
		14'h1a5d: data = 9'o10;
		14'h1a5e: data = 9'o10;
		14'h1a5f: data = 9'o10;
		14'h1a60: data = 9'o21;
		14'h1a61: data = 9'o21;
		14'h1a62: data = 9'o31;
		14'h1a63: data = 9'o142;
		14'h1a64: data = 9'o152;
		14'h1a65: data = 9'o152;
		14'h1a66: data = 9'o152;
		14'h1a67: data = 9'o152;
		14'h1a68: data = 9'o52;
		14'h1a69: data = 9'o52;
		14'h1a6a: data = 9'o52;
		14'h1a6b: data = 9'o273;
		14'h1a6c: data = 9'o272;
		14'h1a6d: data = 9'o172;
		14'h1a6e: data = 9'o172;
		14'h1a6f: data = 9'o172;
		14'h1a70: data = 9'o172;
		14'h1a71: data = 9'o172;
		14'h1a72: data = 9'o172;
		14'h1a73: data = 9'o172;
		14'h1a74: data = 9'o172;
		14'h1a75: data = 9'o172;
		14'h1a76: data = 9'o172;
		14'h1a77: data = 9'o172;
		14'h1a78: data = 9'o172;
		14'h1a79: data = 9'o172;
		14'h1a7a: data = 9'o172;
		14'h1a7b: data = 9'o172;
		14'h1a7c: data = 9'o172;
		14'h1a7d: data = 9'o172;
		14'h1a7e: data = 9'o172;
		14'h1a7f: data = 9'o172;
		14'h1a80: data = 9'o172;
		14'h1a81: data = 9'o272;
		14'h1a82: data = 9'o372;
		14'h1a83: data = 9'o573;
		14'h1a84: data = 9'o773;
		14'h1a85: data = 9'o762;
		14'h1a86: data = 9'o0;
		14'h1a87: data = 9'o0;
		14'h1a88: data = 9'o0;
		14'h1a89: data = 9'o0;
		14'h1a8a: data = 9'o0;
		14'h1a8b: data = 9'o0;
		14'h1a8c: data = 9'o0;
		14'h1a8d: data = 9'o0;
		14'h1a8e: data = 9'o0;
		14'h1a8f: data = 9'o0;
		14'h1a90: data = 9'o0;
		14'h1a91: data = 9'o0;
		14'h1a92: data = 9'o0;
		14'h1a93: data = 9'o0;
		14'h1a94: data = 9'o0;
		14'h1a95: data = 9'o0;
		14'h1a96: data = 9'o0;
		14'h1a97: data = 9'o651;
		14'h1a98: data = 9'o662;
		14'h1a99: data = 9'o773;
		14'h1a9a: data = 9'o573;
		14'h1a9b: data = 9'o372;
		14'h1a9c: data = 9'o272;
		14'h1a9d: data = 9'o172;
		14'h1a9e: data = 9'o172;
		14'h1a9f: data = 9'o172;
		14'h1aa0: data = 9'o172;
		14'h1aa1: data = 9'o172;
		14'h1aa2: data = 9'o172;
		14'h1aa3: data = 9'o172;
		14'h1aa4: data = 9'o172;
		14'h1aa5: data = 9'o172;
		14'h1aa6: data = 9'o172;
		14'h1aa7: data = 9'o172;
		14'h1aa8: data = 9'o172;
		14'h1aa9: data = 9'o172;
		14'h1aaa: data = 9'o172;
		14'h1aab: data = 9'o172;
		14'h1aac: data = 9'o172;
		14'h1aad: data = 9'o172;
		14'h1aae: data = 9'o172;
		14'h1aaf: data = 9'o172;
		14'h1ab0: data = 9'o172;
		14'h1ab1: data = 9'o273;
		14'h1ab2: data = 9'o273;
		14'h1ab3: data = 9'o52;
		14'h1ab4: data = 9'o52;
		14'h1ab5: data = 9'o52;
		14'h1ab6: data = 9'o152;
		14'h1ab7: data = 9'o152;
		14'h1ab8: data = 9'o152;
		14'h1ab9: data = 9'o142;
		14'h1aba: data = 9'o31;
		14'h1abb: data = 9'o21;
		14'h1abc: data = 9'o10;
		14'h1abd: data = 9'o10;
		14'h1abe: data = 9'o11;
		14'h1abf: data = 9'o10;
		14'h1ac0: data = 9'o10;
		14'h1ac1: data = 9'o10;
		14'h1ac2: data = 9'o10;
		14'h1ac3: data = 9'o10;
		14'h1ac4: data = 9'o10;
		14'h1ac5: data = 9'o10;
		14'h1ac6: data = 9'o21;
		14'h1ac7: data = 9'o21;
		14'h1ac8: data = 9'o142;
		14'h1ac9: data = 9'o152;
		14'h1aca: data = 9'o152;
		14'h1acb: data = 9'o152;
		14'h1acc: data = 9'o152;
		14'h1acd: data = 9'o52;
		14'h1ace: data = 9'o52;
		14'h1acf: data = 9'o273;
		14'h1ad0: data = 9'o272;
		14'h1ad1: data = 9'o172;
		14'h1ad2: data = 9'o172;
		14'h1ad3: data = 9'o172;
		14'h1ad4: data = 9'o172;
		14'h1ad5: data = 9'o172;
		14'h1ad6: data = 9'o172;
		14'h1ad7: data = 9'o172;
		14'h1ad8: data = 9'o172;
		14'h1ad9: data = 9'o172;
		14'h1ada: data = 9'o172;
		14'h1adb: data = 9'o172;
		14'h1adc: data = 9'o172;
		14'h1add: data = 9'o172;
		14'h1ade: data = 9'o172;
		14'h1adf: data = 9'o172;
		14'h1ae0: data = 9'o172;
		14'h1ae1: data = 9'o172;
		14'h1ae2: data = 9'o172;
		14'h1ae3: data = 9'o172;
		14'h1ae4: data = 9'o172;
		14'h1ae5: data = 9'o272;
		14'h1ae6: data = 9'o272;
		14'h1ae7: data = 9'o573;
		14'h1ae8: data = 9'o773;
		14'h1ae9: data = 9'o762;
		14'h1aea: data = 9'o0;
		14'h1aeb: data = 9'o0;
		14'h1aec: data = 9'o0;
		14'h1aed: data = 9'o0;
		14'h1aee: data = 9'o0;
		14'h1aef: data = 9'o0;
		14'h1af0: data = 9'o0;
		14'h1af1: data = 9'o0;
		14'h1af2: data = 9'o0;
		14'h1af3: data = 9'o0;
		14'h1af4: data = 9'o0;
		14'h1af5: data = 9'o0;
		14'h1af6: data = 9'o0;
		14'h1af7: data = 9'o0;
		14'h1af8: data = 9'o0;
		14'h1af9: data = 9'o0;
		14'h1afa: data = 9'o0;
		14'h1afb: data = 9'o651;
		14'h1afc: data = 9'o662;
		14'h1afd: data = 9'o773;
		14'h1afe: data = 9'o573;
		14'h1aff: data = 9'o272;
		14'h1b00: data = 9'o272;
		14'h1b01: data = 9'o172;
		14'h1b02: data = 9'o172;
		14'h1b03: data = 9'o172;
		14'h1b04: data = 9'o172;
		14'h1b05: data = 9'o172;
		14'h1b06: data = 9'o172;
		14'h1b07: data = 9'o172;
		14'h1b08: data = 9'o172;
		14'h1b09: data = 9'o172;
		14'h1b0a: data = 9'o172;
		14'h1b0b: data = 9'o172;
		14'h1b0c: data = 9'o172;
		14'h1b0d: data = 9'o172;
		14'h1b0e: data = 9'o172;
		14'h1b0f: data = 9'o172;
		14'h1b10: data = 9'o172;
		14'h1b11: data = 9'o172;
		14'h1b12: data = 9'o172;
		14'h1b13: data = 9'o172;
		14'h1b14: data = 9'o172;
		14'h1b15: data = 9'o273;
		14'h1b16: data = 9'o273;
		14'h1b17: data = 9'o52;
		14'h1b18: data = 9'o52;
		14'h1b19: data = 9'o152;
		14'h1b1a: data = 9'o52;
		14'h1b1b: data = 9'o152;
		14'h1b1c: data = 9'o142;
		14'h1b1d: data = 9'o21;
		14'h1b1e: data = 9'o11;
		14'h1b1f: data = 9'o11;
		14'h1b20: data = 9'o10;
		14'h1b21: data = 9'o10;
		14'h1b22: data = 9'o10;
		14'h1b23: data = 9'o10;
		14'h1b24: data = 9'o10;
		14'h1b25: data = 9'o10;
		14'h1b26: data = 9'o10;
		14'h1b27: data = 9'o10;
		14'h1b28: data = 9'o10;
		14'h1b29: data = 9'o10;
		14'h1b2a: data = 9'o10;
		14'h1b2b: data = 9'o10;
		14'h1b2c: data = 9'o31;
		14'h1b2d: data = 9'o142;
		14'h1b2e: data = 9'o152;
		14'h1b2f: data = 9'o152;
		14'h1b30: data = 9'o152;
		14'h1b31: data = 9'o52;
		14'h1b32: data = 9'o52;
		14'h1b33: data = 9'o273;
		14'h1b34: data = 9'o272;
		14'h1b35: data = 9'o172;
		14'h1b36: data = 9'o172;
		14'h1b37: data = 9'o172;
		14'h1b38: data = 9'o172;
		14'h1b39: data = 9'o172;
		14'h1b3a: data = 9'o172;
		14'h1b3b: data = 9'o172;
		14'h1b3c: data = 9'o172;
		14'h1b3d: data = 9'o172;
		14'h1b3e: data = 9'o172;
		14'h1b3f: data = 9'o172;
		14'h1b40: data = 9'o172;
		14'h1b41: data = 9'o172;
		14'h1b42: data = 9'o172;
		14'h1b43: data = 9'o172;
		14'h1b44: data = 9'o172;
		14'h1b45: data = 9'o172;
		14'h1b46: data = 9'o172;
		14'h1b47: data = 9'o172;
		14'h1b48: data = 9'o172;
		14'h1b49: data = 9'o272;
		14'h1b4a: data = 9'o272;
		14'h1b4b: data = 9'o573;
		14'h1b4c: data = 9'o773;
		14'h1b4d: data = 9'o762;
		14'h1b4e: data = 9'o0;
		14'h1b4f: data = 9'o0;
		14'h1b50: data = 9'o0;
		14'h1b51: data = 9'o0;
		14'h1b52: data = 9'o0;
		14'h1b53: data = 9'o0;
		14'h1b54: data = 9'o0;
		14'h1b55: data = 9'o0;
		14'h1b56: data = 9'o0;
		14'h1b57: data = 9'o0;
		14'h1b58: data = 9'o0;
		14'h1b59: data = 9'o0;
		14'h1b5a: data = 9'o0;
		14'h1b5b: data = 9'o0;
		14'h1b5c: data = 9'o0;
		14'h1b5d: data = 9'o0;
		14'h1b5e: data = 9'o0;
		14'h1b5f: data = 9'o651;
		14'h1b60: data = 9'o662;
		14'h1b61: data = 9'o773;
		14'h1b62: data = 9'o473;
		14'h1b63: data = 9'o272;
		14'h1b64: data = 9'o272;
		14'h1b65: data = 9'o172;
		14'h1b66: data = 9'o272;
		14'h1b67: data = 9'o172;
		14'h1b68: data = 9'o172;
		14'h1b69: data = 9'o172;
		14'h1b6a: data = 9'o172;
		14'h1b6b: data = 9'o172;
		14'h1b6c: data = 9'o172;
		14'h1b6d: data = 9'o172;
		14'h1b6e: data = 9'o172;
		14'h1b6f: data = 9'o172;
		14'h1b70: data = 9'o172;
		14'h1b71: data = 9'o172;
		14'h1b72: data = 9'o172;
		14'h1b73: data = 9'o172;
		14'h1b74: data = 9'o172;
		14'h1b75: data = 9'o172;
		14'h1b76: data = 9'o172;
		14'h1b77: data = 9'o172;
		14'h1b78: data = 9'o172;
		14'h1b79: data = 9'o273;
		14'h1b7a: data = 9'o273;
		14'h1b7b: data = 9'o52;
		14'h1b7c: data = 9'o52;
		14'h1b7d: data = 9'o152;
		14'h1b7e: data = 9'o152;
		14'h1b7f: data = 9'o142;
		14'h1b80: data = 9'o31;
		14'h1b81: data = 9'o10;
		14'h1b82: data = 9'o10;
		14'h1b83: data = 9'o11;
		14'h1b84: data = 9'o10;
		14'h1b85: data = 9'o10;
		14'h1b86: data = 9'o10;
		14'h1b87: data = 9'o10;
		14'h1b88: data = 9'o10;
		14'h1b89: data = 9'o10;
		14'h1b8a: data = 9'o10;
		14'h1b8b: data = 9'o10;
		14'h1b8c: data = 9'o10;
		14'h1b8d: data = 9'o10;
		14'h1b8e: data = 9'o11;
		14'h1b8f: data = 9'o10;
		14'h1b90: data = 9'o10;
		14'h1b91: data = 9'o31;
		14'h1b92: data = 9'o142;
		14'h1b93: data = 9'o152;
		14'h1b94: data = 9'o152;
		14'h1b95: data = 9'o152;
		14'h1b96: data = 9'o52;
		14'h1b97: data = 9'o273;
		14'h1b98: data = 9'o272;
		14'h1b99: data = 9'o172;
		14'h1b9a: data = 9'o172;
		14'h1b9b: data = 9'o172;
		14'h1b9c: data = 9'o172;
		14'h1b9d: data = 9'o172;
		14'h1b9e: data = 9'o172;
		14'h1b9f: data = 9'o172;
		14'h1ba0: data = 9'o172;
		14'h1ba1: data = 9'o172;
		14'h1ba2: data = 9'o172;
		14'h1ba3: data = 9'o172;
		14'h1ba4: data = 9'o172;
		14'h1ba5: data = 9'o172;
		14'h1ba6: data = 9'o172;
		14'h1ba7: data = 9'o172;
		14'h1ba8: data = 9'o172;
		14'h1ba9: data = 9'o172;
		14'h1baa: data = 9'o172;
		14'h1bab: data = 9'o172;
		14'h1bac: data = 9'o172;
		14'h1bad: data = 9'o272;
		14'h1bae: data = 9'o272;
		14'h1baf: data = 9'o473;
		14'h1bb0: data = 9'o773;
		14'h1bb1: data = 9'o762;
		14'h1bb2: data = 9'o0;
		14'h1bb3: data = 9'o0;
		14'h1bb4: data = 9'o0;
		14'h1bb5: data = 9'o0;
		14'h1bb6: data = 9'o0;
		14'h1bb7: data = 9'o0;
		14'h1bb8: data = 9'o0;
		14'h1bb9: data = 9'o0;
		14'h1bba: data = 9'o0;
		14'h1bbb: data = 9'o0;
		14'h1bbc: data = 9'o0;
		14'h1bbd: data = 9'o0;
		14'h1bbe: data = 9'o0;
		14'h1bbf: data = 9'o0;
		14'h1bc0: data = 9'o0;
		14'h1bc1: data = 9'o0;
		14'h1bc2: data = 9'o0;
		14'h1bc3: data = 9'o651;
		14'h1bc4: data = 9'o662;
		14'h1bc5: data = 9'o773;
		14'h1bc6: data = 9'o473;
		14'h1bc7: data = 9'o272;
		14'h1bc8: data = 9'o272;
		14'h1bc9: data = 9'o272;
		14'h1bca: data = 9'o272;
		14'h1bcb: data = 9'o172;
		14'h1bcc: data = 9'o172;
		14'h1bcd: data = 9'o172;
		14'h1bce: data = 9'o172;
		14'h1bcf: data = 9'o172;
		14'h1bd0: data = 9'o172;
		14'h1bd1: data = 9'o172;
		14'h1bd2: data = 9'o172;
		14'h1bd3: data = 9'o172;
		14'h1bd4: data = 9'o172;
		14'h1bd5: data = 9'o172;
		14'h1bd6: data = 9'o172;
		14'h1bd7: data = 9'o172;
		14'h1bd8: data = 9'o172;
		14'h1bd9: data = 9'o172;
		14'h1bda: data = 9'o172;
		14'h1bdb: data = 9'o172;
		14'h1bdc: data = 9'o172;
		14'h1bdd: data = 9'o273;
		14'h1bde: data = 9'o273;
		14'h1bdf: data = 9'o52;
		14'h1be0: data = 9'o52;
		14'h1be1: data = 9'o152;
		14'h1be2: data = 9'o152;
		14'h1be3: data = 9'o31;
		14'h1be4: data = 9'o21;
		14'h1be5: data = 9'o10;
		14'h1be6: data = 9'o10;
		14'h1be7: data = 9'o10;
		14'h1be8: data = 9'o10;
		14'h1be9: data = 9'o10;
		14'h1bea: data = 9'o10;
		14'h1beb: data = 9'o10;
		14'h1bec: data = 9'o10;
		14'h1bed: data = 9'o10;
		14'h1bee: data = 9'o10;
		14'h1bef: data = 9'o10;
		14'h1bf0: data = 9'o11;
		14'h1bf1: data = 9'o11;
		14'h1bf2: data = 9'o10;
		14'h1bf3: data = 9'o10;
		14'h1bf4: data = 9'o10;
		14'h1bf5: data = 9'o21;
		14'h1bf6: data = 9'o32;
		14'h1bf7: data = 9'o152;
		14'h1bf8: data = 9'o152;
		14'h1bf9: data = 9'o152;
		14'h1bfa: data = 9'o52;
		14'h1bfb: data = 9'o273;
		14'h1bfc: data = 9'o272;
		14'h1bfd: data = 9'o172;
		14'h1bfe: data = 9'o172;
		14'h1bff: data = 9'o172;
		14'h1c00: data = 9'o272;
		14'h1c01: data = 9'o272;
		14'h1c02: data = 9'o172;
		14'h1c03: data = 9'o172;
		14'h1c04: data = 9'o172;
		14'h1c05: data = 9'o172;
		14'h1c06: data = 9'o172;
		14'h1c07: data = 9'o172;
		14'h1c08: data = 9'o172;
		14'h1c09: data = 9'o172;
		14'h1c0a: data = 9'o172;
		14'h1c0b: data = 9'o172;
		14'h1c0c: data = 9'o172;
		14'h1c0d: data = 9'o172;
		14'h1c0e: data = 9'o172;
		14'h1c0f: data = 9'o172;
		14'h1c10: data = 9'o172;
		14'h1c11: data = 9'o272;
		14'h1c12: data = 9'o272;
		14'h1c13: data = 9'o473;
		14'h1c14: data = 9'o773;
		14'h1c15: data = 9'o762;
		14'h1c16: data = 9'o0;
		14'h1c17: data = 9'o0;
		14'h1c18: data = 9'o0;
		14'h1c19: data = 9'o0;
		14'h1c1a: data = 9'o0;
		14'h1c1b: data = 9'o0;
		14'h1c1c: data = 9'o0;
		14'h1c1d: data = 9'o0;
		14'h1c1e: data = 9'o0;
		14'h1c1f: data = 9'o0;
		14'h1c20: data = 9'o0;
		14'h1c21: data = 9'o0;
		14'h1c22: data = 9'o0;
		14'h1c23: data = 9'o0;
		14'h1c24: data = 9'o0;
		14'h1c25: data = 9'o0;
		14'h1c26: data = 9'o0;
		14'h1c27: data = 9'o651;
		14'h1c28: data = 9'o662;
		14'h1c29: data = 9'o773;
		14'h1c2a: data = 9'o473;
		14'h1c2b: data = 9'o272;
		14'h1c2c: data = 9'o272;
		14'h1c2d: data = 9'o272;
		14'h1c2e: data = 9'o272;
		14'h1c2f: data = 9'o272;
		14'h1c30: data = 9'o172;
		14'h1c31: data = 9'o172;
		14'h1c32: data = 9'o172;
		14'h1c33: data = 9'o172;
		14'h1c34: data = 9'o172;
		14'h1c35: data = 9'o172;
		14'h1c36: data = 9'o172;
		14'h1c37: data = 9'o172;
		14'h1c38: data = 9'o172;
		14'h1c39: data = 9'o172;
		14'h1c3a: data = 9'o172;
		14'h1c3b: data = 9'o172;
		14'h1c3c: data = 9'o172;
		14'h1c3d: data = 9'o172;
		14'h1c3e: data = 9'o172;
		14'h1c3f: data = 9'o172;
		14'h1c40: data = 9'o172;
		14'h1c41: data = 9'o273;
		14'h1c42: data = 9'o173;
		14'h1c43: data = 9'o52;
		14'h1c44: data = 9'o52;
		14'h1c45: data = 9'o152;
		14'h1c46: data = 9'o142;
		14'h1c47: data = 9'o21;
		14'h1c48: data = 9'o10;
		14'h1c49: data = 9'o10;
		14'h1c4a: data = 9'o10;
		14'h1c4b: data = 9'o10;
		14'h1c4c: data = 9'o10;
		14'h1c4d: data = 9'o10;
		14'h1c4e: data = 9'o10;
		14'h1c4f: data = 9'o10;
		14'h1c50: data = 9'o10;
		14'h1c51: data = 9'o10;
		14'h1c52: data = 9'o10;
		14'h1c53: data = 9'o10;
		14'h1c54: data = 9'o10;
		14'h1c55: data = 9'o10;
		14'h1c56: data = 9'o10;
		14'h1c57: data = 9'o10;
		14'h1c58: data = 9'o10;
		14'h1c59: data = 9'o10;
		14'h1c5a: data = 9'o21;
		14'h1c5b: data = 9'o142;
		14'h1c5c: data = 9'o152;
		14'h1c5d: data = 9'o52;
		14'h1c5e: data = 9'o52;
		14'h1c5f: data = 9'o273;
		14'h1c60: data = 9'o272;
		14'h1c61: data = 9'o172;
		14'h1c62: data = 9'o172;
		14'h1c63: data = 9'o172;
		14'h1c64: data = 9'o172;
		14'h1c65: data = 9'o272;
		14'h1c66: data = 9'o172;
		14'h1c67: data = 9'o172;
		14'h1c68: data = 9'o172;
		14'h1c69: data = 9'o172;
		14'h1c6a: data = 9'o172;
		14'h1c6b: data = 9'o172;
		14'h1c6c: data = 9'o172;
		14'h1c6d: data = 9'o172;
		14'h1c6e: data = 9'o172;
		14'h1c6f: data = 9'o172;
		14'h1c70: data = 9'o172;
		14'h1c71: data = 9'o172;
		14'h1c72: data = 9'o172;
		14'h1c73: data = 9'o172;
		14'h1c74: data = 9'o172;
		14'h1c75: data = 9'o172;
		14'h1c76: data = 9'o272;
		14'h1c77: data = 9'o373;
		14'h1c78: data = 9'o773;
		14'h1c79: data = 9'o763;
		14'h1c7a: data = 9'o0;
		14'h1c7b: data = 9'o0;
		14'h1c7c: data = 9'o0;
		14'h1c7d: data = 9'o0;
		14'h1c7e: data = 9'o0;
		14'h1c7f: data = 9'o0;
		14'h1c80: data = 9'o0;
		14'h1c81: data = 9'o0;
		14'h1c82: data = 9'o0;
		14'h1c83: data = 9'o0;
		14'h1c84: data = 9'o0;
		14'h1c85: data = 9'o0;
		14'h1c86: data = 9'o0;
		14'h1c87: data = 9'o0;
		14'h1c88: data = 9'o0;
		14'h1c89: data = 9'o0;
		14'h1c8a: data = 9'o0;
		14'h1c8b: data = 9'o641;
		14'h1c8c: data = 9'o662;
		14'h1c8d: data = 9'o773;
		14'h1c8e: data = 9'o372;
		14'h1c8f: data = 9'o272;
		14'h1c90: data = 9'o172;
		14'h1c91: data = 9'o172;
		14'h1c92: data = 9'o272;
		14'h1c93: data = 9'o272;
		14'h1c94: data = 9'o172;
		14'h1c95: data = 9'o172;
		14'h1c96: data = 9'o172;
		14'h1c97: data = 9'o172;
		14'h1c98: data = 9'o172;
		14'h1c99: data = 9'o172;
		14'h1c9a: data = 9'o172;
		14'h1c9b: data = 9'o172;
		14'h1c9c: data = 9'o172;
		14'h1c9d: data = 9'o172;
		14'h1c9e: data = 9'o172;
		14'h1c9f: data = 9'o172;
		14'h1ca0: data = 9'o172;
		14'h1ca1: data = 9'o172;
		14'h1ca2: data = 9'o172;
		14'h1ca3: data = 9'o172;
		14'h1ca4: data = 9'o172;
		14'h1ca5: data = 9'o173;
		14'h1ca6: data = 9'o173;
		14'h1ca7: data = 9'o52;
		14'h1ca8: data = 9'o152;
		14'h1ca9: data = 9'o152;
		14'h1caa: data = 9'o31;
		14'h1cab: data = 9'o21;
		14'h1cac: data = 9'o10;
		14'h1cad: data = 9'o10;
		14'h1cae: data = 9'o10;
		14'h1caf: data = 9'o10;
		14'h1cb0: data = 9'o10;
		14'h1cb1: data = 9'o10;
		14'h1cb2: data = 9'o10;
		14'h1cb3: data = 9'o10;
		14'h1cb4: data = 9'o10;
		14'h1cb5: data = 9'o10;
		14'h1cb6: data = 9'o10;
		14'h1cb7: data = 9'o10;
		14'h1cb8: data = 9'o10;
		14'h1cb9: data = 9'o10;
		14'h1cba: data = 9'o10;
		14'h1cbb: data = 9'o10;
		14'h1cbc: data = 9'o10;
		14'h1cbd: data = 9'o10;
		14'h1cbe: data = 9'o21;
		14'h1cbf: data = 9'o31;
		14'h1cc0: data = 9'o252;
		14'h1cc1: data = 9'o152;
		14'h1cc2: data = 9'o152;
		14'h1cc3: data = 9'o172;
		14'h1cc4: data = 9'o173;
		14'h1cc5: data = 9'o172;
		14'h1cc6: data = 9'o172;
		14'h1cc7: data = 9'o172;
		14'h1cc8: data = 9'o172;
		14'h1cc9: data = 9'o272;
		14'h1cca: data = 9'o172;
		14'h1ccb: data = 9'o172;
		14'h1ccc: data = 9'o172;
		14'h1ccd: data = 9'o172;
		14'h1cce: data = 9'o172;
		14'h1ccf: data = 9'o172;
		14'h1cd0: data = 9'o172;
		14'h1cd1: data = 9'o172;
		14'h1cd2: data = 9'o172;
		14'h1cd3: data = 9'o172;
		14'h1cd4: data = 9'o172;
		14'h1cd5: data = 9'o172;
		14'h1cd6: data = 9'o172;
		14'h1cd7: data = 9'o172;
		14'h1cd8: data = 9'o172;
		14'h1cd9: data = 9'o172;
		14'h1cda: data = 9'o272;
		14'h1cdb: data = 9'o373;
		14'h1cdc: data = 9'o673;
		14'h1cdd: data = 9'o763;
		14'h1cde: data = 9'o0;
		14'h1cdf: data = 9'o0;
		14'h1ce0: data = 9'o0;
		14'h1ce1: data = 9'o0;
		14'h1ce2: data = 9'o0;
		14'h1ce3: data = 9'o0;
		14'h1ce4: data = 9'o0;
		14'h1ce5: data = 9'o0;
		14'h1ce6: data = 9'o0;
		14'h1ce7: data = 9'o0;
		14'h1ce8: data = 9'o0;
		14'h1ce9: data = 9'o0;
		14'h1cea: data = 9'o0;
		14'h1ceb: data = 9'o0;
		14'h1cec: data = 9'o0;
		14'h1ced: data = 9'o0;
		14'h1cee: data = 9'o0;
		14'h1cef: data = 9'o641;
		14'h1cf0: data = 9'o662;
		14'h1cf1: data = 9'o773;
		14'h1cf2: data = 9'o372;
		14'h1cf3: data = 9'o272;
		14'h1cf4: data = 9'o172;
		14'h1cf5: data = 9'o172;
		14'h1cf6: data = 9'o272;
		14'h1cf7: data = 9'o272;
		14'h1cf8: data = 9'o172;
		14'h1cf9: data = 9'o172;
		14'h1cfa: data = 9'o172;
		14'h1cfb: data = 9'o172;
		14'h1cfc: data = 9'o172;
		14'h1cfd: data = 9'o172;
		14'h1cfe: data = 9'o172;
		14'h1cff: data = 9'o172;
		14'h1d00: data = 9'o172;
		14'h1d01: data = 9'o172;
		14'h1d02: data = 9'o172;
		14'h1d03: data = 9'o172;
		14'h1d04: data = 9'o172;
		14'h1d05: data = 9'o172;
		14'h1d06: data = 9'o172;
		14'h1d07: data = 9'o172;
		14'h1d08: data = 9'o172;
		14'h1d09: data = 9'o273;
		14'h1d0a: data = 9'o273;
		14'h1d0b: data = 9'o52;
		14'h1d0c: data = 9'o152;
		14'h1d0d: data = 9'o142;
		14'h1d0e: data = 9'o21;
		14'h1d0f: data = 9'o10;
		14'h1d10: data = 9'o10;
		14'h1d11: data = 9'o10;
		14'h1d12: data = 9'o10;
		14'h1d13: data = 9'o10;
		14'h1d14: data = 9'o10;
		14'h1d15: data = 9'o10;
		14'h1d16: data = 9'o10;
		14'h1d17: data = 9'o10;
		14'h1d18: data = 9'o10;
		14'h1d19: data = 9'o10;
		14'h1d1a: data = 9'o10;
		14'h1d1b: data = 9'o10;
		14'h1d1c: data = 9'o10;
		14'h1d1d: data = 9'o10;
		14'h1d1e: data = 9'o10;
		14'h1d1f: data = 9'o10;
		14'h1d20: data = 9'o10;
		14'h1d21: data = 9'o11;
		14'h1d22: data = 9'o11;
		14'h1d23: data = 9'o21;
		14'h1d24: data = 9'o142;
		14'h1d25: data = 9'o152;
		14'h1d26: data = 9'o152;
		14'h1d27: data = 9'o173;
		14'h1d28: data = 9'o273;
		14'h1d29: data = 9'o172;
		14'h1d2a: data = 9'o172;
		14'h1d2b: data = 9'o172;
		14'h1d2c: data = 9'o172;
		14'h1d2d: data = 9'o172;
		14'h1d2e: data = 9'o172;
		14'h1d2f: data = 9'o172;
		14'h1d30: data = 9'o172;
		14'h1d31: data = 9'o172;
		14'h1d32: data = 9'o172;
		14'h1d33: data = 9'o172;
		14'h1d34: data = 9'o172;
		14'h1d35: data = 9'o172;
		14'h1d36: data = 9'o172;
		14'h1d37: data = 9'o172;
		14'h1d38: data = 9'o172;
		14'h1d39: data = 9'o172;
		14'h1d3a: data = 9'o172;
		14'h1d3b: data = 9'o172;
		14'h1d3c: data = 9'o172;
		14'h1d3d: data = 9'o172;
		14'h1d3e: data = 9'o172;
		14'h1d3f: data = 9'o372;
		14'h1d40: data = 9'o673;
		14'h1d41: data = 9'o673;
		14'h1d42: data = 9'o0;
		14'h1d43: data = 9'o0;
		14'h1d44: data = 9'o0;
		14'h1d45: data = 9'o0;
		14'h1d46: data = 9'o0;
		14'h1d47: data = 9'o0;
		14'h1d48: data = 9'o0;
		14'h1d49: data = 9'o0;
		14'h1d4a: data = 9'o0;
		14'h1d4b: data = 9'o0;
		14'h1d4c: data = 9'o0;
		14'h1d4d: data = 9'o0;
		14'h1d4e: data = 9'o0;
		14'h1d4f: data = 9'o0;
		14'h1d50: data = 9'o0;
		14'h1d51: data = 9'o0;
		14'h1d52: data = 9'o0;
		14'h1d53: data = 9'o541;
		14'h1d54: data = 9'o662;
		14'h1d55: data = 9'o673;
		14'h1d56: data = 9'o372;
		14'h1d57: data = 9'o272;
		14'h1d58: data = 9'o172;
		14'h1d59: data = 9'o172;
		14'h1d5a: data = 9'o272;
		14'h1d5b: data = 9'o272;
		14'h1d5c: data = 9'o172;
		14'h1d5d: data = 9'o172;
		14'h1d5e: data = 9'o172;
		14'h1d5f: data = 9'o172;
		14'h1d60: data = 9'o172;
		14'h1d61: data = 9'o172;
		14'h1d62: data = 9'o172;
		14'h1d63: data = 9'o172;
		14'h1d64: data = 9'o172;
		14'h1d65: data = 9'o272;
		14'h1d66: data = 9'o272;
		14'h1d67: data = 9'o272;
		14'h1d68: data = 9'o272;
		14'h1d69: data = 9'o172;
		14'h1d6a: data = 9'o172;
		14'h1d6b: data = 9'o172;
		14'h1d6c: data = 9'o172;
		14'h1d6d: data = 9'o272;
		14'h1d6e: data = 9'o273;
		14'h1d6f: data = 9'o152;
		14'h1d70: data = 9'o152;
		14'h1d71: data = 9'o142;
		14'h1d72: data = 9'o21;
		14'h1d73: data = 9'o10;
		14'h1d74: data = 9'o10;
		14'h1d75: data = 9'o10;
		14'h1d76: data = 9'o10;
		14'h1d77: data = 9'o10;
		14'h1d78: data = 9'o10;
		14'h1d79: data = 9'o10;
		14'h1d7a: data = 9'o10;
		14'h1d7b: data = 9'o10;
		14'h1d7c: data = 9'o10;
		14'h1d7d: data = 9'o10;
		14'h1d7e: data = 9'o10;
		14'h1d7f: data = 9'o10;
		14'h1d80: data = 9'o10;
		14'h1d81: data = 9'o10;
		14'h1d82: data = 9'o10;
		14'h1d83: data = 9'o10;
		14'h1d84: data = 9'o10;
		14'h1d85: data = 9'o10;
		14'h1d86: data = 9'o10;
		14'h1d87: data = 9'o21;
		14'h1d88: data = 9'o142;
		14'h1d89: data = 9'o152;
		14'h1d8a: data = 9'o52;
		14'h1d8b: data = 9'o172;
		14'h1d8c: data = 9'o173;
		14'h1d8d: data = 9'o172;
		14'h1d8e: data = 9'o172;
		14'h1d8f: data = 9'o172;
		14'h1d90: data = 9'o172;
		14'h1d91: data = 9'o172;
		14'h1d92: data = 9'o172;
		14'h1d93: data = 9'o172;
		14'h1d94: data = 9'o172;
		14'h1d95: data = 9'o172;
		14'h1d96: data = 9'o172;
		14'h1d97: data = 9'o172;
		14'h1d98: data = 9'o172;
		14'h1d99: data = 9'o172;
		14'h1d9a: data = 9'o172;
		14'h1d9b: data = 9'o172;
		14'h1d9c: data = 9'o172;
		14'h1d9d: data = 9'o172;
		14'h1d9e: data = 9'o172;
		14'h1d9f: data = 9'o172;
		14'h1da0: data = 9'o172;
		14'h1da1: data = 9'o272;
		14'h1da2: data = 9'o272;
		14'h1da3: data = 9'o372;
		14'h1da4: data = 9'o673;
		14'h1da5: data = 9'o673;
		14'h1da6: data = 9'o0;
		14'h1da7: data = 9'o0;
		14'h1da8: data = 9'o0;
		14'h1da9: data = 9'o0;
		14'h1daa: data = 9'o0;
		14'h1dab: data = 9'o0;
		14'h1dac: data = 9'o0;
		14'h1dad: data = 9'o0;
		14'h1dae: data = 9'o0;
		14'h1daf: data = 9'o0;
		14'h1db0: data = 9'o0;
		14'h1db1: data = 9'o0;
		14'h1db2: data = 9'o0;
		14'h1db3: data = 9'o0;
		14'h1db4: data = 9'o0;
		14'h1db5: data = 9'o0;
		14'h1db6: data = 9'o0;
		14'h1db7: data = 9'o551;
		14'h1db8: data = 9'o662;
		14'h1db9: data = 9'o673;
		14'h1dba: data = 9'o272;
		14'h1dbb: data = 9'o172;
		14'h1dbc: data = 9'o172;
		14'h1dbd: data = 9'o172;
		14'h1dbe: data = 9'o272;
		14'h1dbf: data = 9'o272;
		14'h1dc0: data = 9'o172;
		14'h1dc1: data = 9'o172;
		14'h1dc2: data = 9'o172;
		14'h1dc3: data = 9'o272;
		14'h1dc4: data = 9'o172;
		14'h1dc5: data = 9'o172;
		14'h1dc6: data = 9'o172;
		14'h1dc7: data = 9'o172;
		14'h1dc8: data = 9'o272;
		14'h1dc9: data = 9'o272;
		14'h1dca: data = 9'o272;
		14'h1dcb: data = 9'o272;
		14'h1dcc: data = 9'o272;
		14'h1dcd: data = 9'o272;
		14'h1dce: data = 9'o272;
		14'h1dcf: data = 9'o272;
		14'h1dd0: data = 9'o172;
		14'h1dd1: data = 9'o272;
		14'h1dd2: data = 9'o272;
		14'h1dd3: data = 9'o52;
		14'h1dd4: data = 9'o152;
		14'h1dd5: data = 9'o142;
		14'h1dd6: data = 9'o10;
		14'h1dd7: data = 9'o10;
		14'h1dd8: data = 9'o10;
		14'h1dd9: data = 9'o10;
		14'h1dda: data = 9'o10;
		14'h1ddb: data = 9'o10;
		14'h1ddc: data = 9'o10;
		14'h1ddd: data = 9'o10;
		14'h1dde: data = 9'o10;
		14'h1ddf: data = 9'o10;
		14'h1de0: data = 9'o10;
		14'h1de1: data = 9'o10;
		14'h1de2: data = 9'o10;
		14'h1de3: data = 9'o10;
		14'h1de4: data = 9'o10;
		14'h1de5: data = 9'o10;
		14'h1de6: data = 9'o10;
		14'h1de7: data = 9'o10;
		14'h1de8: data = 9'o10;
		14'h1de9: data = 9'o10;
		14'h1dea: data = 9'o11;
		14'h1deb: data = 9'o21;
		14'h1dec: data = 9'o142;
		14'h1ded: data = 9'o152;
		14'h1dee: data = 9'o152;
		14'h1def: data = 9'o273;
		14'h1df0: data = 9'o273;
		14'h1df1: data = 9'o172;
		14'h1df2: data = 9'o172;
		14'h1df3: data = 9'o172;
		14'h1df4: data = 9'o272;
		14'h1df5: data = 9'o172;
		14'h1df6: data = 9'o272;
		14'h1df7: data = 9'o272;
		14'h1df8: data = 9'o272;
		14'h1df9: data = 9'o272;
		14'h1dfa: data = 9'o272;
		14'h1dfb: data = 9'o272;
		14'h1dfc: data = 9'o272;
		14'h1dfd: data = 9'o272;
		14'h1dfe: data = 9'o272;
		14'h1dff: data = 9'o272;
		14'h1e00: data = 9'o272;
		14'h1e01: data = 9'o272;
		14'h1e02: data = 9'o272;
		14'h1e03: data = 9'o272;
		14'h1e04: data = 9'o272;
		14'h1e05: data = 9'o272;
		14'h1e06: data = 9'o272;
		14'h1e07: data = 9'o272;
		14'h1e08: data = 9'o673;
		14'h1e09: data = 9'o662;
		14'h1e0a: data = 9'o0;
		14'h1e0b: data = 9'o0;
		14'h1e0c: data = 9'o0;
		14'h1e0d: data = 9'o0;
		14'h1e0e: data = 9'o0;
		14'h1e0f: data = 9'o0;
		14'h1e10: data = 9'o0;
		14'h1e11: data = 9'o0;
		14'h1e12: data = 9'o0;
		14'h1e13: data = 9'o0;
		14'h1e14: data = 9'o0;
		14'h1e15: data = 9'o0;
		14'h1e16: data = 9'o0;
		14'h1e17: data = 9'o0;
		14'h1e18: data = 9'o0;
		14'h1e19: data = 9'o0;
		14'h1e1a: data = 9'o0;
		14'h1e1b: data = 9'o551;
		14'h1e1c: data = 9'o662;
		14'h1e1d: data = 9'o673;
		14'h1e1e: data = 9'o372;
		14'h1e1f: data = 9'o172;
		14'h1e20: data = 9'o172;
		14'h1e21: data = 9'o172;
		14'h1e22: data = 9'o172;
		14'h1e23: data = 9'o172;
		14'h1e24: data = 9'o172;
		14'h1e25: data = 9'o172;
		14'h1e26: data = 9'o172;
		14'h1e27: data = 9'o172;
		14'h1e28: data = 9'o172;
		14'h1e29: data = 9'o172;
		14'h1e2a: data = 9'o172;
		14'h1e2b: data = 9'o172;
		14'h1e2c: data = 9'o172;
		14'h1e2d: data = 9'o172;
		14'h1e2e: data = 9'o172;
		14'h1e2f: data = 9'o172;
		14'h1e30: data = 9'o172;
		14'h1e31: data = 9'o172;
		14'h1e32: data = 9'o172;
		14'h1e33: data = 9'o172;
		14'h1e34: data = 9'o172;
		14'h1e35: data = 9'o272;
		14'h1e36: data = 9'o273;
		14'h1e37: data = 9'o52;
		14'h1e38: data = 9'o52;
		14'h1e39: data = 9'o42;
		14'h1e3a: data = 9'o10;
		14'h1e3b: data = 9'o10;
		14'h1e3c: data = 9'o10;
		14'h1e3d: data = 9'o10;
		14'h1e3e: data = 9'o10;
		14'h1e3f: data = 9'o10;
		14'h1e40: data = 9'o10;
		14'h1e41: data = 9'o10;
		14'h1e42: data = 9'o10;
		14'h1e43: data = 9'o10;
		14'h1e44: data = 9'o10;
		14'h1e45: data = 9'o10;
		14'h1e46: data = 9'o10;
		14'h1e47: data = 9'o10;
		14'h1e48: data = 9'o10;
		14'h1e49: data = 9'o10;
		14'h1e4a: data = 9'o10;
		14'h1e4b: data = 9'o10;
		14'h1e4c: data = 9'o10;
		14'h1e4d: data = 9'o10;
		14'h1e4e: data = 9'o21;
		14'h1e4f: data = 9'o21;
		14'h1e50: data = 9'o31;
		14'h1e51: data = 9'o152;
		14'h1e52: data = 9'o152;
		14'h1e53: data = 9'o272;
		14'h1e54: data = 9'o273;
		14'h1e55: data = 9'o172;
		14'h1e56: data = 9'o172;
		14'h1e57: data = 9'o172;
		14'h1e58: data = 9'o172;
		14'h1e59: data = 9'o172;
		14'h1e5a: data = 9'o172;
		14'h1e5b: data = 9'o172;
		14'h1e5c: data = 9'o172;
		14'h1e5d: data = 9'o172;
		14'h1e5e: data = 9'o172;
		14'h1e5f: data = 9'o172;
		14'h1e60: data = 9'o172;
		14'h1e61: data = 9'o172;
		14'h1e62: data = 9'o172;
		14'h1e63: data = 9'o172;
		14'h1e64: data = 9'o172;
		14'h1e65: data = 9'o172;
		14'h1e66: data = 9'o172;
		14'h1e67: data = 9'o172;
		14'h1e68: data = 9'o172;
		14'h1e69: data = 9'o172;
		14'h1e6a: data = 9'o272;
		14'h1e6b: data = 9'o272;
		14'h1e6c: data = 9'o573;
		14'h1e6d: data = 9'o673;
		14'h1e6e: data = 9'o0;
		14'h1e6f: data = 9'o0;
		14'h1e70: data = 9'o0;
		14'h1e71: data = 9'o0;
		14'h1e72: data = 9'o0;
		14'h1e73: data = 9'o0;
		14'h1e74: data = 9'o0;
		14'h1e75: data = 9'o0;
		14'h1e76: data = 9'o0;
		14'h1e77: data = 9'o0;
		14'h1e78: data = 9'o0;
		14'h1e79: data = 9'o0;
		14'h1e7a: data = 9'o0;
		14'h1e7b: data = 9'o0;
		14'h1e7c: data = 9'o0;
		14'h1e7d: data = 9'o0;
		14'h1e7e: data = 9'o0;
		14'h1e7f: data = 9'o551;
		14'h1e80: data = 9'o662;
		14'h1e81: data = 9'o573;
		14'h1e82: data = 9'o372;
		14'h1e83: data = 9'o272;
		14'h1e84: data = 9'o272;
		14'h1e85: data = 9'o272;
		14'h1e86: data = 9'o272;
		14'h1e87: data = 9'o272;
		14'h1e88: data = 9'o272;
		14'h1e89: data = 9'o272;
		14'h1e8a: data = 9'o272;
		14'h1e8b: data = 9'o272;
		14'h1e8c: data = 9'o272;
		14'h1e8d: data = 9'o272;
		14'h1e8e: data = 9'o272;
		14'h1e8f: data = 9'o272;
		14'h1e90: data = 9'o272;
		14'h1e91: data = 9'o272;
		14'h1e92: data = 9'o272;
		14'h1e93: data = 9'o272;
		14'h1e94: data = 9'o272;
		14'h1e95: data = 9'o272;
		14'h1e96: data = 9'o272;
		14'h1e97: data = 9'o272;
		14'h1e98: data = 9'o272;
		14'h1e99: data = 9'o272;
		14'h1e9a: data = 9'o272;
		14'h1e9b: data = 9'o152;
		14'h1e9c: data = 9'o152;
		14'h1e9d: data = 9'o41;
		14'h1e9e: data = 9'o10;
		14'h1e9f: data = 9'o10;
		14'h1ea0: data = 9'o10;
		14'h1ea1: data = 9'o10;
		14'h1ea2: data = 9'o10;
		14'h1ea3: data = 9'o10;
		14'h1ea4: data = 9'o10;
		14'h1ea5: data = 9'o10;
		14'h1ea6: data = 9'o10;
		14'h1ea7: data = 9'o10;
		14'h1ea8: data = 9'o10;
		14'h1ea9: data = 9'o10;
		14'h1eaa: data = 9'o10;
		14'h1eab: data = 9'o10;
		14'h1eac: data = 9'o10;
		14'h1ead: data = 9'o10;
		14'h1eae: data = 9'o10;
		14'h1eaf: data = 9'o10;
		14'h1eb0: data = 9'o10;
		14'h1eb1: data = 9'o10;
		14'h1eb2: data = 9'o10;
		14'h1eb3: data = 9'o20;
		14'h1eb4: data = 9'o31;
		14'h1eb5: data = 9'o152;
		14'h1eb6: data = 9'o152;
		14'h1eb7: data = 9'o272;
		14'h1eb8: data = 9'o273;
		14'h1eb9: data = 9'o272;
		14'h1eba: data = 9'o272;
		14'h1ebb: data = 9'o272;
		14'h1ebc: data = 9'o272;
		14'h1ebd: data = 9'o272;
		14'h1ebe: data = 9'o272;
		14'h1ebf: data = 9'o272;
		14'h1ec0: data = 9'o272;
		14'h1ec1: data = 9'o272;
		14'h1ec2: data = 9'o272;
		14'h1ec3: data = 9'o272;
		14'h1ec4: data = 9'o272;
		14'h1ec5: data = 9'o272;
		14'h1ec6: data = 9'o272;
		14'h1ec7: data = 9'o272;
		14'h1ec8: data = 9'o272;
		14'h1ec9: data = 9'o272;
		14'h1eca: data = 9'o272;
		14'h1ecb: data = 9'o272;
		14'h1ecc: data = 9'o272;
		14'h1ecd: data = 9'o272;
		14'h1ece: data = 9'o272;
		14'h1ecf: data = 9'o372;
		14'h1ed0: data = 9'o573;
		14'h1ed1: data = 9'o673;
		14'h1ed2: data = 9'o0;
		14'h1ed3: data = 9'o0;
		14'h1ed4: data = 9'o0;
		14'h1ed5: data = 9'o0;
		14'h1ed6: data = 9'o0;
		14'h1ed7: data = 9'o0;
		14'h1ed8: data = 9'o0;
		14'h1ed9: data = 9'o0;
		14'h1eda: data = 9'o0;
		14'h1edb: data = 9'o0;
		14'h1edc: data = 9'o0;
		14'h1edd: data = 9'o0;
		14'h1ede: data = 9'o0;
		14'h1edf: data = 9'o0;
		14'h1ee0: data = 9'o0;
		14'h1ee1: data = 9'o0;
		14'h1ee2: data = 9'o0;
		14'h1ee3: data = 9'o551;
		14'h1ee4: data = 9'o662;
		14'h1ee5: data = 9'o673;
		14'h1ee6: data = 9'o372;
		14'h1ee7: data = 9'o372;
		14'h1ee8: data = 9'o372;
		14'h1ee9: data = 9'o272;
		14'h1eea: data = 9'o372;
		14'h1eeb: data = 9'o372;
		14'h1eec: data = 9'o272;
		14'h1eed: data = 9'o272;
		14'h1eee: data = 9'o372;
		14'h1eef: data = 9'o372;
		14'h1ef0: data = 9'o372;
		14'h1ef1: data = 9'o372;
		14'h1ef2: data = 9'o372;
		14'h1ef3: data = 9'o372;
		14'h1ef4: data = 9'o372;
		14'h1ef5: data = 9'o372;
		14'h1ef6: data = 9'o372;
		14'h1ef7: data = 9'o372;
		14'h1ef8: data = 9'o372;
		14'h1ef9: data = 9'o372;
		14'h1efa: data = 9'o372;
		14'h1efb: data = 9'o372;
		14'h1efc: data = 9'o372;
		14'h1efd: data = 9'o372;
		14'h1efe: data = 9'o362;
		14'h1eff: data = 9'o252;
		14'h1f00: data = 9'o252;
		14'h1f01: data = 9'o142;
		14'h1f02: data = 9'o10;
		14'h1f03: data = 9'o10;
		14'h1f04: data = 9'o10;
		14'h1f05: data = 9'o10;
		14'h1f06: data = 9'o10;
		14'h1f07: data = 9'o10;
		14'h1f08: data = 9'o10;
		14'h1f09: data = 9'o10;
		14'h1f0a: data = 9'o10;
		14'h1f0b: data = 9'o10;
		14'h1f0c: data = 9'o10;
		14'h1f0d: data = 9'o10;
		14'h1f0e: data = 9'o10;
		14'h1f0f: data = 9'o10;
		14'h1f10: data = 9'o10;
		14'h1f11: data = 9'o10;
		14'h1f12: data = 9'o10;
		14'h1f13: data = 9'o10;
		14'h1f14: data = 9'o10;
		14'h1f15: data = 9'o10;
		14'h1f16: data = 9'o11;
		14'h1f17: data = 9'o21;
		14'h1f18: data = 9'o131;
		14'h1f19: data = 9'o242;
		14'h1f1a: data = 9'o252;
		14'h1f1b: data = 9'o362;
		14'h1f1c: data = 9'o372;
		14'h1f1d: data = 9'o372;
		14'h1f1e: data = 9'o372;
		14'h1f1f: data = 9'o372;
		14'h1f20: data = 9'o372;
		14'h1f21: data = 9'o372;
		14'h1f22: data = 9'o372;
		14'h1f23: data = 9'o372;
		14'h1f24: data = 9'o372;
		14'h1f25: data = 9'o372;
		14'h1f26: data = 9'o372;
		14'h1f27: data = 9'o372;
		14'h1f28: data = 9'o372;
		14'h1f29: data = 9'o372;
		14'h1f2a: data = 9'o372;
		14'h1f2b: data = 9'o372;
		14'h1f2c: data = 9'o372;
		14'h1f2d: data = 9'o372;
		14'h1f2e: data = 9'o372;
		14'h1f2f: data = 9'o372;
		14'h1f30: data = 9'o372;
		14'h1f31: data = 9'o372;
		14'h1f32: data = 9'o372;
		14'h1f33: data = 9'o372;
		14'h1f34: data = 9'o573;
		14'h1f35: data = 9'o662;
		14'h1f36: data = 9'o0;
		14'h1f37: data = 9'o0;
		14'h1f38: data = 9'o0;
		14'h1f39: data = 9'o0;
		14'h1f3a: data = 9'o0;
		14'h1f3b: data = 9'o0;
		14'h1f3c: data = 9'o0;
		14'h1f3d: data = 9'o0;
		14'h1f3e: data = 9'o0;
		14'h1f3f: data = 9'o0;
		14'h1f40: data = 9'o0;
		14'h1f41: data = 9'o0;
		14'h1f42: data = 9'o0;
		14'h1f43: data = 9'o0;
		14'h1f44: data = 9'o0;
		14'h1f45: data = 9'o0;
		14'h1f46: data = 9'o0;
		14'h1f47: data = 9'o551;
		14'h1f48: data = 9'o662;
		14'h1f49: data = 9'o773;
		14'h1f4a: data = 9'o573;
		14'h1f4b: data = 9'o573;
		14'h1f4c: data = 9'o573;
		14'h1f4d: data = 9'o573;
		14'h1f4e: data = 9'o573;
		14'h1f4f: data = 9'o573;
		14'h1f50: data = 9'o573;
		14'h1f51: data = 9'o573;
		14'h1f52: data = 9'o573;
		14'h1f53: data = 9'o573;
		14'h1f54: data = 9'o573;
		14'h1f55: data = 9'o573;
		14'h1f56: data = 9'o573;
		14'h1f57: data = 9'o573;
		14'h1f58: data = 9'o573;
		14'h1f59: data = 9'o573;
		14'h1f5a: data = 9'o573;
		14'h1f5b: data = 9'o573;
		14'h1f5c: data = 9'o573;
		14'h1f5d: data = 9'o573;
		14'h1f5e: data = 9'o573;
		14'h1f5f: data = 9'o573;
		14'h1f60: data = 9'o573;
		14'h1f61: data = 9'o573;
		14'h1f62: data = 9'o673;
		14'h1f63: data = 9'o573;
		14'h1f64: data = 9'o673;
		14'h1f65: data = 9'o673;
		14'h1f66: data = 9'o673;
		14'h1f67: data = 9'o673;
		14'h1f68: data = 9'o673;
		14'h1f69: data = 9'o673;
		14'h1f6a: data = 9'o663;
		14'h1f6b: data = 9'o663;
		14'h1f6c: data = 9'o663;
		14'h1f6d: data = 9'o663;
		14'h1f6e: data = 9'o663;
		14'h1f6f: data = 9'o663;
		14'h1f70: data = 9'o663;
		14'h1f71: data = 9'o663;
		14'h1f72: data = 9'o663;
		14'h1f73: data = 9'o663;
		14'h1f74: data = 9'o663;
		14'h1f75: data = 9'o663;
		14'h1f76: data = 9'o663;
		14'h1f77: data = 9'o663;
		14'h1f78: data = 9'o663;
		14'h1f79: data = 9'o673;
		14'h1f7a: data = 9'o673;
		14'h1f7b: data = 9'o673;
		14'h1f7c: data = 9'o673;
		14'h1f7d: data = 9'o673;
		14'h1f7e: data = 9'o573;
		14'h1f7f: data = 9'o673;
		14'h1f80: data = 9'o573;
		14'h1f81: data = 9'o573;
		14'h1f82: data = 9'o573;
		14'h1f83: data = 9'o573;
		14'h1f84: data = 9'o573;
		14'h1f85: data = 9'o573;
		14'h1f86: data = 9'o573;
		14'h1f87: data = 9'o573;
		14'h1f88: data = 9'o573;
		14'h1f89: data = 9'o573;
		14'h1f8a: data = 9'o573;
		14'h1f8b: data = 9'o573;
		14'h1f8c: data = 9'o573;
		14'h1f8d: data = 9'o573;
		14'h1f8e: data = 9'o573;
		14'h1f8f: data = 9'o573;
		14'h1f90: data = 9'o573;
		14'h1f91: data = 9'o573;
		14'h1f92: data = 9'o573;
		14'h1f93: data = 9'o573;
		14'h1f94: data = 9'o573;
		14'h1f95: data = 9'o573;
		14'h1f96: data = 9'o573;
		14'h1f97: data = 9'o673;
		14'h1f98: data = 9'o773;
		14'h1f99: data = 9'o773;
		14'h1f9a: data = 9'o0;
		14'h1f9b: data = 9'o0;
		14'h1f9c: data = 9'o0;
		14'h1f9d: data = 9'o0;
		14'h1f9e: data = 9'o0;
		14'h1f9f: data = 9'o0;
		14'h1fa0: data = 9'o0;
		14'h1fa1: data = 9'o0;
		14'h1fa2: data = 9'o0;
		14'h1fa3: data = 9'o0;
		14'h1fa4: data = 9'o0;
		14'h1fa5: data = 9'o0;
		14'h1fa6: data = 9'o0;
		14'h1fa7: data = 9'o0;
		14'h1fa8: data = 9'o0;
		14'h1fa9: data = 9'o0;
		14'h1faa: data = 9'o0;
		14'h1fab: data = 9'o651;
		14'h1fac: data = 9'o762;
		14'h1fad: data = 9'o773;
		14'h1fae: data = 9'o773;
		14'h1faf: data = 9'o773;
		14'h1fb0: data = 9'o773;
		14'h1fb1: data = 9'o773;
		14'h1fb2: data = 9'o773;
		14'h1fb3: data = 9'o773;
		14'h1fb4: data = 9'o773;
		14'h1fb5: data = 9'o773;
		14'h1fb6: data = 9'o773;
		14'h1fb7: data = 9'o773;
		14'h1fb8: data = 9'o773;
		14'h1fb9: data = 9'o773;
		14'h1fba: data = 9'o773;
		14'h1fbb: data = 9'o773;
		14'h1fbc: data = 9'o773;
		14'h1fbd: data = 9'o773;
		14'h1fbe: data = 9'o773;
		14'h1fbf: data = 9'o773;
		14'h1fc0: data = 9'o773;
		14'h1fc1: data = 9'o773;
		14'h1fc2: data = 9'o773;
		14'h1fc3: data = 9'o773;
		14'h1fc4: data = 9'o773;
		14'h1fc5: data = 9'o773;
		14'h1fc6: data = 9'o773;
		14'h1fc7: data = 9'o773;
		14'h1fc8: data = 9'o773;
		14'h1fc9: data = 9'o773;
		14'h1fca: data = 9'o773;
		14'h1fcb: data = 9'o773;
		14'h1fcc: data = 9'o773;
		14'h1fcd: data = 9'o773;
		14'h1fce: data = 9'o773;
		14'h1fcf: data = 9'o773;
		14'h1fd0: data = 9'o773;
		14'h1fd1: data = 9'o773;
		14'h1fd2: data = 9'o773;
		14'h1fd3: data = 9'o773;
		14'h1fd4: data = 9'o773;
		14'h1fd5: data = 9'o773;
		14'h1fd6: data = 9'o773;
		14'h1fd7: data = 9'o773;
		14'h1fd8: data = 9'o773;
		14'h1fd9: data = 9'o773;
		14'h1fda: data = 9'o773;
		14'h1fdb: data = 9'o773;
		14'h1fdc: data = 9'o773;
		14'h1fdd: data = 9'o773;
		14'h1fde: data = 9'o773;
		14'h1fdf: data = 9'o773;
		14'h1fe0: data = 9'o773;
		14'h1fe1: data = 9'o773;
		14'h1fe2: data = 9'o773;
		14'h1fe3: data = 9'o773;
		14'h1fe4: data = 9'o773;
		14'h1fe5: data = 9'o773;
		14'h1fe6: data = 9'o773;
		14'h1fe7: data = 9'o773;
		14'h1fe8: data = 9'o773;
		14'h1fe9: data = 9'o773;
		14'h1fea: data = 9'o773;
		14'h1feb: data = 9'o773;
		14'h1fec: data = 9'o773;
		14'h1fed: data = 9'o773;
		14'h1fee: data = 9'o773;
		14'h1fef: data = 9'o773;
		14'h1ff0: data = 9'o773;
		14'h1ff1: data = 9'o773;
		14'h1ff2: data = 9'o773;
		14'h1ff3: data = 9'o773;
		14'h1ff4: data = 9'o773;
		14'h1ff5: data = 9'o773;
		14'h1ff6: data = 9'o773;
		14'h1ff7: data = 9'o773;
		14'h1ff8: data = 9'o773;
		14'h1ff9: data = 9'o773;
		14'h1ffa: data = 9'o773;
		14'h1ffb: data = 9'o773;
		14'h1ffc: data = 9'o773;
		14'h1ffd: data = 9'o763;
		14'h1ffe: data = 9'o0;
		14'h1fff: data = 9'o0;
		14'h2000: data = 9'o0;
		14'h2001: data = 9'o0;
		14'h2002: data = 9'o0;
		14'h2003: data = 9'o0;
		14'h2004: data = 9'o0;
		14'h2005: data = 9'o0;
		14'h2006: data = 9'o0;
		14'h2007: data = 9'o0;
		14'h2008: data = 9'o0;
		14'h2009: data = 9'o0;
		14'h200a: data = 9'o0;
		14'h200b: data = 9'o0;
		14'h200c: data = 9'o0;
		14'h200d: data = 9'o0;
		14'h200e: data = 9'o0;
		14'h200f: data = 9'o651;
		14'h2010: data = 9'o762;
		14'h2011: data = 9'o773;
		14'h2012: data = 9'o773;
		14'h2013: data = 9'o773;
		14'h2014: data = 9'o773;
		14'h2015: data = 9'o773;
		14'h2016: data = 9'o773;
		14'h2017: data = 9'o773;
		14'h2018: data = 9'o773;
		14'h2019: data = 9'o773;
		14'h201a: data = 9'o773;
		14'h201b: data = 9'o773;
		14'h201c: data = 9'o773;
		14'h201d: data = 9'o773;
		14'h201e: data = 9'o773;
		14'h201f: data = 9'o773;
		14'h2020: data = 9'o773;
		14'h2021: data = 9'o773;
		14'h2022: data = 9'o773;
		14'h2023: data = 9'o773;
		14'h2024: data = 9'o773;
		14'h2025: data = 9'o773;
		14'h2026: data = 9'o773;
		14'h2027: data = 9'o773;
		14'h2028: data = 9'o773;
		14'h2029: data = 9'o773;
		14'h202a: data = 9'o773;
		14'h202b: data = 9'o773;
		14'h202c: data = 9'o773;
		14'h202d: data = 9'o773;
		14'h202e: data = 9'o773;
		14'h202f: data = 9'o773;
		14'h2030: data = 9'o773;
		14'h2031: data = 9'o773;
		14'h2032: data = 9'o773;
		14'h2033: data = 9'o773;
		14'h2034: data = 9'o773;
		14'h2035: data = 9'o773;
		14'h2036: data = 9'o773;
		14'h2037: data = 9'o773;
		14'h2038: data = 9'o773;
		14'h2039: data = 9'o773;
		14'h203a: data = 9'o773;
		14'h203b: data = 9'o773;
		14'h203c: data = 9'o773;
		14'h203d: data = 9'o773;
		14'h203e: data = 9'o773;
		14'h203f: data = 9'o773;
		14'h2040: data = 9'o773;
		14'h2041: data = 9'o773;
		14'h2042: data = 9'o773;
		14'h2043: data = 9'o773;
		14'h2044: data = 9'o773;
		14'h2045: data = 9'o773;
		14'h2046: data = 9'o773;
		14'h2047: data = 9'o773;
		14'h2048: data = 9'o773;
		14'h2049: data = 9'o773;
		14'h204a: data = 9'o773;
		14'h204b: data = 9'o773;
		14'h204c: data = 9'o773;
		14'h204d: data = 9'o773;
		14'h204e: data = 9'o773;
		14'h204f: data = 9'o773;
		14'h2050: data = 9'o773;
		14'h2051: data = 9'o773;
		14'h2052: data = 9'o773;
		14'h2053: data = 9'o773;
		14'h2054: data = 9'o773;
		14'h2055: data = 9'o773;
		14'h2056: data = 9'o773;
		14'h2057: data = 9'o773;
		14'h2058: data = 9'o773;
		14'h2059: data = 9'o773;
		14'h205a: data = 9'o773;
		14'h205b: data = 9'o773;
		14'h205c: data = 9'o773;
		14'h205d: data = 9'o773;
		14'h205e: data = 9'o773;
		14'h205f: data = 9'o773;
		14'h2060: data = 9'o773;
		14'h2061: data = 9'o762;
		14'h2062: data = 9'o0;
		14'h2063: data = 9'o0;
		14'h2064: data = 9'o0;
		14'h2065: data = 9'o0;
		14'h2066: data = 9'o0;
		14'h2067: data = 9'o0;
		14'h2068: data = 9'o0;
		14'h2069: data = 9'o0;
		14'h206a: data = 9'o0;
		14'h206b: data = 9'o0;
		14'h206c: data = 9'o0;
		14'h206d: data = 9'o0;
		14'h206e: data = 9'o0;
		14'h206f: data = 9'o0;
		14'h2070: data = 9'o0;
		14'h2071: data = 9'o0;
		14'h2072: data = 9'o0;
		14'h2073: data = 9'o651;
		14'h2074: data = 9'o662;
		14'h2075: data = 9'o773;
		14'h2076: data = 9'o773;
		14'h2077: data = 9'o773;
		14'h2078: data = 9'o773;
		14'h2079: data = 9'o773;
		14'h207a: data = 9'o773;
		14'h207b: data = 9'o773;
		14'h207c: data = 9'o773;
		14'h207d: data = 9'o773;
		14'h207e: data = 9'o773;
		14'h207f: data = 9'o773;
		14'h2080: data = 9'o773;
		14'h2081: data = 9'o773;
		14'h2082: data = 9'o773;
		14'h2083: data = 9'o773;
		14'h2084: data = 9'o773;
		14'h2085: data = 9'o773;
		14'h2086: data = 9'o773;
		14'h2087: data = 9'o773;
		14'h2088: data = 9'o773;
		14'h2089: data = 9'o773;
		14'h208a: data = 9'o773;
		14'h208b: data = 9'o773;
		14'h208c: data = 9'o773;
		14'h208d: data = 9'o773;
		14'h208e: data = 9'o773;
		14'h208f: data = 9'o773;
		14'h2090: data = 9'o773;
		14'h2091: data = 9'o773;
		14'h2092: data = 9'o773;
		14'h2093: data = 9'o773;
		14'h2094: data = 9'o773;
		14'h2095: data = 9'o773;
		14'h2096: data = 9'o773;
		14'h2097: data = 9'o773;
		14'h2098: data = 9'o773;
		14'h2099: data = 9'o773;
		14'h209a: data = 9'o773;
		14'h209b: data = 9'o773;
		14'h209c: data = 9'o773;
		14'h209d: data = 9'o773;
		14'h209e: data = 9'o773;
		14'h209f: data = 9'o773;
		14'h20a0: data = 9'o773;
		14'h20a1: data = 9'o773;
		14'h20a2: data = 9'o773;
		14'h20a3: data = 9'o773;
		14'h20a4: data = 9'o773;
		14'h20a5: data = 9'o773;
		14'h20a6: data = 9'o773;
		14'h20a7: data = 9'o773;
		14'h20a8: data = 9'o773;
		14'h20a9: data = 9'o773;
		14'h20aa: data = 9'o773;
		14'h20ab: data = 9'o773;
		14'h20ac: data = 9'o773;
		14'h20ad: data = 9'o773;
		14'h20ae: data = 9'o773;
		14'h20af: data = 9'o773;
		14'h20b0: data = 9'o773;
		14'h20b1: data = 9'o773;
		14'h20b2: data = 9'o773;
		14'h20b3: data = 9'o773;
		14'h20b4: data = 9'o773;
		14'h20b5: data = 9'o773;
		14'h20b6: data = 9'o773;
		14'h20b7: data = 9'o773;
		14'h20b8: data = 9'o773;
		14'h20b9: data = 9'o773;
		14'h20ba: data = 9'o773;
		14'h20bb: data = 9'o773;
		14'h20bc: data = 9'o773;
		14'h20bd: data = 9'o773;
		14'h20be: data = 9'o773;
		14'h20bf: data = 9'o773;
		14'h20c0: data = 9'o773;
		14'h20c1: data = 9'o773;
		14'h20c2: data = 9'o773;
		14'h20c3: data = 9'o773;
		14'h20c4: data = 9'o773;
		14'h20c5: data = 9'o762;
		14'h20c6: data = 9'o0;
		14'h20c7: data = 9'o0;
		14'h20c8: data = 9'o0;
		14'h20c9: data = 9'o0;
		14'h20ca: data = 9'o0;
		14'h20cb: data = 9'o0;
		14'h20cc: data = 9'o0;
		14'h20cd: data = 9'o0;
		14'h20ce: data = 9'o0;
		14'h20cf: data = 9'o0;
		14'h20d0: data = 9'o0;
		14'h20d1: data = 9'o0;
		14'h20d2: data = 9'o0;
		14'h20d3: data = 9'o0;
		14'h20d4: data = 9'o0;
		14'h20d5: data = 9'o0;
		14'h20d6: data = 9'o0;
		14'h20d7: data = 9'o651;
		14'h20d8: data = 9'o662;
		14'h20d9: data = 9'o773;
		14'h20da: data = 9'o773;
		14'h20db: data = 9'o773;
		14'h20dc: data = 9'o773;
		14'h20dd: data = 9'o773;
		14'h20de: data = 9'o773;
		14'h20df: data = 9'o773;
		14'h20e0: data = 9'o773;
		14'h20e1: data = 9'o773;
		14'h20e2: data = 9'o773;
		14'h20e3: data = 9'o773;
		14'h20e4: data = 9'o773;
		14'h20e5: data = 9'o773;
		14'h20e6: data = 9'o773;
		14'h20e7: data = 9'o773;
		14'h20e8: data = 9'o773;
		14'h20e9: data = 9'o773;
		14'h20ea: data = 9'o773;
		14'h20eb: data = 9'o773;
		14'h20ec: data = 9'o773;
		14'h20ed: data = 9'o773;
		14'h20ee: data = 9'o773;
		14'h20ef: data = 9'o773;
		14'h20f0: data = 9'o773;
		14'h20f1: data = 9'o773;
		14'h20f2: data = 9'o773;
		14'h20f3: data = 9'o773;
		14'h20f4: data = 9'o773;
		14'h20f5: data = 9'o773;
		14'h20f6: data = 9'o773;
		14'h20f7: data = 9'o773;
		14'h20f8: data = 9'o773;
		14'h20f9: data = 9'o773;
		14'h20fa: data = 9'o773;
		14'h20fb: data = 9'o773;
		14'h20fc: data = 9'o773;
		14'h20fd: data = 9'o773;
		14'h20fe: data = 9'o773;
		14'h20ff: data = 9'o773;
		14'h2100: data = 9'o773;
		14'h2101: data = 9'o773;
		14'h2102: data = 9'o773;
		14'h2103: data = 9'o773;
		14'h2104: data = 9'o773;
		14'h2105: data = 9'o773;
		14'h2106: data = 9'o773;
		14'h2107: data = 9'o773;
		14'h2108: data = 9'o773;
		14'h2109: data = 9'o773;
		14'h210a: data = 9'o773;
		14'h210b: data = 9'o773;
		14'h210c: data = 9'o773;
		14'h210d: data = 9'o773;
		14'h210e: data = 9'o773;
		14'h210f: data = 9'o773;
		14'h2110: data = 9'o773;
		14'h2111: data = 9'o773;
		14'h2112: data = 9'o773;
		14'h2113: data = 9'o773;
		14'h2114: data = 9'o773;
		14'h2115: data = 9'o773;
		14'h2116: data = 9'o773;
		14'h2117: data = 9'o773;
		14'h2118: data = 9'o773;
		14'h2119: data = 9'o773;
		14'h211a: data = 9'o773;
		14'h211b: data = 9'o773;
		14'h211c: data = 9'o773;
		14'h211d: data = 9'o773;
		14'h211e: data = 9'o773;
		14'h211f: data = 9'o773;
		14'h2120: data = 9'o773;
		14'h2121: data = 9'o773;
		14'h2122: data = 9'o773;
		14'h2123: data = 9'o773;
		14'h2124: data = 9'o773;
		14'h2125: data = 9'o773;
		14'h2126: data = 9'o773;
		14'h2127: data = 9'o773;
		14'h2128: data = 9'o773;
		14'h2129: data = 9'o662;
		14'h212a: data = 9'o0;
		14'h212b: data = 9'o0;
		14'h212c: data = 9'o0;
		14'h212d: data = 9'o0;
		14'h212e: data = 9'o0;
		14'h212f: data = 9'o0;
		14'h2130: data = 9'o0;
		14'h2131: data = 9'o0;
		14'h2132: data = 9'o0;
		14'h2133: data = 9'o0;
		14'h2134: data = 9'o0;
		14'h2135: data = 9'o0;
		14'h2136: data = 9'o0;
		14'h2137: data = 9'o0;
		14'h2138: data = 9'o0;
		14'h2139: data = 9'o0;
		14'h213a: data = 9'o0;
		14'h213b: data = 9'o551;
		14'h213c: data = 9'o662;
		14'h213d: data = 9'o773;
		14'h213e: data = 9'o773;
		14'h213f: data = 9'o773;
		14'h2140: data = 9'o773;
		14'h2141: data = 9'o773;
		14'h2142: data = 9'o773;
		14'h2143: data = 9'o773;
		14'h2144: data = 9'o773;
		14'h2145: data = 9'o773;
		14'h2146: data = 9'o773;
		14'h2147: data = 9'o773;
		14'h2148: data = 9'o773;
		14'h2149: data = 9'o773;
		14'h214a: data = 9'o773;
		14'h214b: data = 9'o773;
		14'h214c: data = 9'o773;
		14'h214d: data = 9'o773;
		14'h214e: data = 9'o773;
		14'h214f: data = 9'o773;
		14'h2150: data = 9'o773;
		14'h2151: data = 9'o773;
		14'h2152: data = 9'o773;
		14'h2153: data = 9'o773;
		14'h2154: data = 9'o773;
		14'h2155: data = 9'o773;
		14'h2156: data = 9'o773;
		14'h2157: data = 9'o773;
		14'h2158: data = 9'o773;
		14'h2159: data = 9'o773;
		14'h215a: data = 9'o773;
		14'h215b: data = 9'o773;
		14'h215c: data = 9'o773;
		14'h215d: data = 9'o773;
		14'h215e: data = 9'o773;
		14'h215f: data = 9'o773;
		14'h2160: data = 9'o773;
		14'h2161: data = 9'o773;
		14'h2162: data = 9'o773;
		14'h2163: data = 9'o773;
		14'h2164: data = 9'o773;
		14'h2165: data = 9'o773;
		14'h2166: data = 9'o773;
		14'h2167: data = 9'o773;
		14'h2168: data = 9'o773;
		14'h2169: data = 9'o773;
		14'h216a: data = 9'o773;
		14'h216b: data = 9'o773;
		14'h216c: data = 9'o773;
		14'h216d: data = 9'o773;
		14'h216e: data = 9'o773;
		14'h216f: data = 9'o773;
		14'h2170: data = 9'o773;
		14'h2171: data = 9'o773;
		14'h2172: data = 9'o773;
		14'h2173: data = 9'o773;
		14'h2174: data = 9'o773;
		14'h2175: data = 9'o773;
		14'h2176: data = 9'o773;
		14'h2177: data = 9'o773;
		14'h2178: data = 9'o773;
		14'h2179: data = 9'o773;
		14'h217a: data = 9'o773;
		14'h217b: data = 9'o773;
		14'h217c: data = 9'o773;
		14'h217d: data = 9'o773;
		14'h217e: data = 9'o773;
		14'h217f: data = 9'o773;
		14'h2180: data = 9'o773;
		14'h2181: data = 9'o773;
		14'h2182: data = 9'o773;
		14'h2183: data = 9'o773;
		14'h2184: data = 9'o773;
		14'h2185: data = 9'o773;
		14'h2186: data = 9'o773;
		14'h2187: data = 9'o773;
		14'h2188: data = 9'o773;
		14'h2189: data = 9'o773;
		14'h218a: data = 9'o773;
		14'h218b: data = 9'o773;
		14'h218c: data = 9'o773;
		14'h218d: data = 9'o663;
		14'h218e: data = 9'o0;
		14'h218f: data = 9'o0;
		14'h2190: data = 9'o0;
		14'h2191: data = 9'o0;
		14'h2192: data = 9'o0;
		14'h2193: data = 9'o0;
		14'h2194: data = 9'o0;
		14'h2195: data = 9'o0;
		14'h2196: data = 9'o0;
		14'h2197: data = 9'o0;
		14'h2198: data = 9'o0;
		14'h2199: data = 9'o0;
		14'h219a: data = 9'o0;
		14'h219b: data = 9'o0;
		14'h219c: data = 9'o0;
		14'h219d: data = 9'o0;
		14'h219e: data = 9'o0;
		14'h219f: data = 9'o551;
		14'h21a0: data = 9'o662;
		14'h21a1: data = 9'o773;
		14'h21a2: data = 9'o773;
		14'h21a3: data = 9'o773;
		14'h21a4: data = 9'o773;
		14'h21a5: data = 9'o773;
		14'h21a6: data = 9'o773;
		14'h21a7: data = 9'o773;
		14'h21a8: data = 9'o773;
		14'h21a9: data = 9'o773;
		14'h21aa: data = 9'o773;
		14'h21ab: data = 9'o773;
		14'h21ac: data = 9'o773;
		14'h21ad: data = 9'o773;
		14'h21ae: data = 9'o773;
		14'h21af: data = 9'o773;
		14'h21b0: data = 9'o773;
		14'h21b1: data = 9'o773;
		14'h21b2: data = 9'o773;
		14'h21b3: data = 9'o773;
		14'h21b4: data = 9'o773;
		14'h21b5: data = 9'o773;
		14'h21b6: data = 9'o773;
		14'h21b7: data = 9'o773;
		14'h21b8: data = 9'o773;
		14'h21b9: data = 9'o773;
		14'h21ba: data = 9'o773;
		14'h21bb: data = 9'o773;
		14'h21bc: data = 9'o773;
		14'h21bd: data = 9'o773;
		14'h21be: data = 9'o773;
		14'h21bf: data = 9'o773;
		14'h21c0: data = 9'o773;
		14'h21c1: data = 9'o773;
		14'h21c2: data = 9'o773;
		14'h21c3: data = 9'o773;
		14'h21c4: data = 9'o773;
		14'h21c5: data = 9'o773;
		14'h21c6: data = 9'o773;
		14'h21c7: data = 9'o773;
		14'h21c8: data = 9'o773;
		14'h21c9: data = 9'o773;
		14'h21ca: data = 9'o773;
		14'h21cb: data = 9'o773;
		14'h21cc: data = 9'o773;
		14'h21cd: data = 9'o773;
		14'h21ce: data = 9'o773;
		14'h21cf: data = 9'o773;
		14'h21d0: data = 9'o773;
		14'h21d1: data = 9'o773;
		14'h21d2: data = 9'o773;
		14'h21d3: data = 9'o773;
		14'h21d4: data = 9'o773;
		14'h21d5: data = 9'o773;
		14'h21d6: data = 9'o773;
		14'h21d7: data = 9'o773;
		14'h21d8: data = 9'o773;
		14'h21d9: data = 9'o773;
		14'h21da: data = 9'o773;
		14'h21db: data = 9'o773;
		14'h21dc: data = 9'o773;
		14'h21dd: data = 9'o773;
		14'h21de: data = 9'o773;
		14'h21df: data = 9'o773;
		14'h21e0: data = 9'o773;
		14'h21e1: data = 9'o773;
		14'h21e2: data = 9'o773;
		14'h21e3: data = 9'o773;
		14'h21e4: data = 9'o773;
		14'h21e5: data = 9'o773;
		14'h21e6: data = 9'o773;
		14'h21e7: data = 9'o773;
		14'h21e8: data = 9'o773;
		14'h21e9: data = 9'o773;
		14'h21ea: data = 9'o773;
		14'h21eb: data = 9'o773;
		14'h21ec: data = 9'o773;
		14'h21ed: data = 9'o773;
		14'h21ee: data = 9'o773;
		14'h21ef: data = 9'o773;
		14'h21f0: data = 9'o773;
		14'h21f1: data = 9'o663;
		14'h21f2: data = 9'o0;
		14'h21f3: data = 9'o0;
		14'h21f4: data = 9'o0;
		14'h21f5: data = 9'o0;
		14'h21f6: data = 9'o0;
		14'h21f7: data = 9'o0;
		14'h21f8: data = 9'o0;
		14'h21f9: data = 9'o0;
		14'h21fa: data = 9'o0;
		14'h21fb: data = 9'o0;
		14'h21fc: data = 9'o0;
		14'h21fd: data = 9'o0;
		14'h21fe: data = 9'o0;
		14'h21ff: data = 9'o0;
		14'h2200: data = 9'o0;
		14'h2201: data = 9'o0;
		14'h2202: data = 9'o0;
		14'h2203: data = 9'o652;
		14'h2204: data = 9'o662;
		14'h2205: data = 9'o773;
		14'h2206: data = 9'o773;
		14'h2207: data = 9'o773;
		14'h2208: data = 9'o773;
		14'h2209: data = 9'o773;
		14'h220a: data = 9'o773;
		14'h220b: data = 9'o773;
		14'h220c: data = 9'o773;
		14'h220d: data = 9'o773;
		14'h220e: data = 9'o773;
		14'h220f: data = 9'o773;
		14'h2210: data = 9'o773;
		14'h2211: data = 9'o773;
		14'h2212: data = 9'o773;
		14'h2213: data = 9'o773;
		14'h2214: data = 9'o773;
		14'h2215: data = 9'o773;
		14'h2216: data = 9'o773;
		14'h2217: data = 9'o773;
		14'h2218: data = 9'o773;
		14'h2219: data = 9'o773;
		14'h221a: data = 9'o773;
		14'h221b: data = 9'o773;
		14'h221c: data = 9'o773;
		14'h221d: data = 9'o773;
		14'h221e: data = 9'o773;
		14'h221f: data = 9'o773;
		14'h2220: data = 9'o773;
		14'h2221: data = 9'o773;
		14'h2222: data = 9'o773;
		14'h2223: data = 9'o773;
		14'h2224: data = 9'o773;
		14'h2225: data = 9'o773;
		14'h2226: data = 9'o773;
		14'h2227: data = 9'o773;
		14'h2228: data = 9'o773;
		14'h2229: data = 9'o773;
		14'h222a: data = 9'o773;
		14'h222b: data = 9'o773;
		14'h222c: data = 9'o773;
		14'h222d: data = 9'o773;
		14'h222e: data = 9'o773;
		14'h222f: data = 9'o773;
		14'h2230: data = 9'o773;
		14'h2231: data = 9'o773;
		14'h2232: data = 9'o773;
		14'h2233: data = 9'o773;
		14'h2234: data = 9'o773;
		14'h2235: data = 9'o773;
		14'h2236: data = 9'o773;
		14'h2237: data = 9'o773;
		14'h2238: data = 9'o773;
		14'h2239: data = 9'o773;
		14'h223a: data = 9'o773;
		14'h223b: data = 9'o773;
		14'h223c: data = 9'o773;
		14'h223d: data = 9'o773;
		14'h223e: data = 9'o773;
		14'h223f: data = 9'o773;
		14'h2240: data = 9'o773;
		14'h2241: data = 9'o773;
		14'h2242: data = 9'o773;
		14'h2243: data = 9'o773;
		14'h2244: data = 9'o773;
		14'h2245: data = 9'o773;
		14'h2246: data = 9'o773;
		14'h2247: data = 9'o773;
		14'h2248: data = 9'o773;
		14'h2249: data = 9'o773;
		14'h224a: data = 9'o773;
		14'h224b: data = 9'o773;
		14'h224c: data = 9'o773;
		14'h224d: data = 9'o773;
		14'h224e: data = 9'o773;
		14'h224f: data = 9'o773;
		14'h2250: data = 9'o773;
		14'h2251: data = 9'o773;
		14'h2252: data = 9'o773;
		14'h2253: data = 9'o773;
		14'h2254: data = 9'o773;
		14'h2255: data = 9'o763;
		14'h2256: data = 9'o0;
		14'h2257: data = 9'o0;
		14'h2258: data = 9'o0;
		14'h2259: data = 9'o0;
		14'h225a: data = 9'o0;
		14'h225b: data = 9'o0;
		14'h225c: data = 9'o0;
		14'h225d: data = 9'o0;
		14'h225e: data = 9'o0;
		14'h225f: data = 9'o0;
		14'h2260: data = 9'o0;
		14'h2261: data = 9'o0;
		14'h2262: data = 9'o0;
		14'h2263: data = 9'o0;
		14'h2264: data = 9'o0;
		14'h2265: data = 9'o0;
		14'h2266: data = 9'o0;
		14'h2267: data = 9'o641;
		14'h2268: data = 9'o662;
		14'h2269: data = 9'o773;
		14'h226a: data = 9'o773;
		14'h226b: data = 9'o773;
		14'h226c: data = 9'o773;
		14'h226d: data = 9'o773;
		14'h226e: data = 9'o773;
		14'h226f: data = 9'o773;
		14'h2270: data = 9'o773;
		14'h2271: data = 9'o773;
		14'h2272: data = 9'o773;
		14'h2273: data = 9'o773;
		14'h2274: data = 9'o773;
		14'h2275: data = 9'o773;
		14'h2276: data = 9'o773;
		14'h2277: data = 9'o773;
		14'h2278: data = 9'o773;
		14'h2279: data = 9'o773;
		14'h227a: data = 9'o773;
		14'h227b: data = 9'o773;
		14'h227c: data = 9'o773;
		14'h227d: data = 9'o773;
		14'h227e: data = 9'o773;
		14'h227f: data = 9'o773;
		14'h2280: data = 9'o773;
		14'h2281: data = 9'o773;
		14'h2282: data = 9'o773;
		14'h2283: data = 9'o773;
		14'h2284: data = 9'o773;
		14'h2285: data = 9'o773;
		14'h2286: data = 9'o773;
		14'h2287: data = 9'o773;
		14'h2288: data = 9'o773;
		14'h2289: data = 9'o773;
		14'h228a: data = 9'o773;
		14'h228b: data = 9'o773;
		14'h228c: data = 9'o773;
		14'h228d: data = 9'o773;
		14'h228e: data = 9'o773;
		14'h228f: data = 9'o773;
		14'h2290: data = 9'o773;
		14'h2291: data = 9'o773;
		14'h2292: data = 9'o773;
		14'h2293: data = 9'o773;
		14'h2294: data = 9'o773;
		14'h2295: data = 9'o773;
		14'h2296: data = 9'o773;
		14'h2297: data = 9'o773;
		14'h2298: data = 9'o773;
		14'h2299: data = 9'o773;
		14'h229a: data = 9'o773;
		14'h229b: data = 9'o773;
		14'h229c: data = 9'o773;
		14'h229d: data = 9'o773;
		14'h229e: data = 9'o773;
		14'h229f: data = 9'o773;
		14'h22a0: data = 9'o773;
		14'h22a1: data = 9'o773;
		14'h22a2: data = 9'o773;
		14'h22a3: data = 9'o773;
		14'h22a4: data = 9'o773;
		14'h22a5: data = 9'o773;
		14'h22a6: data = 9'o773;
		14'h22a7: data = 9'o773;
		14'h22a8: data = 9'o773;
		14'h22a9: data = 9'o773;
		14'h22aa: data = 9'o773;
		14'h22ab: data = 9'o773;
		14'h22ac: data = 9'o773;
		14'h22ad: data = 9'o773;
		14'h22ae: data = 9'o773;
		14'h22af: data = 9'o773;
		14'h22b0: data = 9'o773;
		14'h22b1: data = 9'o773;
		14'h22b2: data = 9'o773;
		14'h22b3: data = 9'o773;
		14'h22b4: data = 9'o773;
		14'h22b5: data = 9'o773;
		14'h22b6: data = 9'o773;
		14'h22b7: data = 9'o773;
		14'h22b8: data = 9'o773;
		14'h22b9: data = 9'o762;
		14'h22ba: data = 9'o0;
		14'h22bb: data = 9'o0;
		14'h22bc: data = 9'o0;
		14'h22bd: data = 9'o0;
		14'h22be: data = 9'o0;
		14'h22bf: data = 9'o0;
		14'h22c0: data = 9'o0;
		14'h22c1: data = 9'o0;
		14'h22c2: data = 9'o0;
		14'h22c3: data = 9'o0;
		14'h22c4: data = 9'o0;
		14'h22c5: data = 9'o0;
		14'h22c6: data = 9'o0;
		14'h22c7: data = 9'o0;
		14'h22c8: data = 9'o0;
		14'h22c9: data = 9'o0;
		14'h22ca: data = 9'o0;
		14'h22cb: data = 9'o651;
		14'h22cc: data = 9'o651;
		14'h22cd: data = 9'o651;
		14'h22ce: data = 9'o551;
		14'h22cf: data = 9'o551;
		14'h22d0: data = 9'o551;
		14'h22d1: data = 9'o551;
		14'h22d2: data = 9'o551;
		14'h22d3: data = 9'o652;
		14'h22d4: data = 9'o551;
		14'h22d5: data = 9'o652;
		14'h22d6: data = 9'o651;
		14'h22d7: data = 9'o651;
		14'h22d8: data = 9'o651;
		14'h22d9: data = 9'o651;
		14'h22da: data = 9'o651;
		14'h22db: data = 9'o652;
		14'h22dc: data = 9'o551;
		14'h22dd: data = 9'o652;
		14'h22de: data = 9'o652;
		14'h22df: data = 9'o551;
		14'h22e0: data = 9'o652;
		14'h22e1: data = 9'o652;
		14'h22e2: data = 9'o651;
		14'h22e3: data = 9'o651;
		14'h22e4: data = 9'o651;
		14'h22e5: data = 9'o652;
		14'h22e6: data = 9'o652;
		14'h22e7: data = 9'o651;
		14'h22e8: data = 9'o651;
		14'h22e9: data = 9'o651;
		14'h22ea: data = 9'o651;
		14'h22eb: data = 9'o652;
		14'h22ec: data = 9'o652;
		14'h22ed: data = 9'o652;
		14'h22ee: data = 9'o652;
		14'h22ef: data = 9'o651;
		14'h22f0: data = 9'o652;
		14'h22f1: data = 9'o652;
		14'h22f2: data = 9'o551;
		14'h22f3: data = 9'o652;
		14'h22f4: data = 9'o652;
		14'h22f5: data = 9'o551;
		14'h22f6: data = 9'o652;
		14'h22f7: data = 9'o652;
		14'h22f8: data = 9'o652;
		14'h22f9: data = 9'o551;
		14'h22fa: data = 9'o651;
		14'h22fb: data = 9'o651;
		14'h22fc: data = 9'o652;
		14'h22fd: data = 9'o651;
		14'h22fe: data = 9'o551;
		14'h22ff: data = 9'o651;
		14'h2300: data = 9'o551;
		14'h2301: data = 9'o551;
		14'h2302: data = 9'o651;
		14'h2303: data = 9'o541;
		14'h2304: data = 9'o651;
		14'h2305: data = 9'o652;
		14'h2306: data = 9'o651;
		14'h2307: data = 9'o652;
		14'h2308: data = 9'o652;
		14'h2309: data = 9'o541;
		14'h230a: data = 9'o551;
		14'h230b: data = 9'o652;
		14'h230c: data = 9'o652;
		14'h230d: data = 9'o651;
		14'h230e: data = 9'o652;
		14'h230f: data = 9'o652;
		14'h2310: data = 9'o551;
		14'h2311: data = 9'o652;
		14'h2312: data = 9'o652;
		14'h2313: data = 9'o551;
		14'h2314: data = 9'o652;
		14'h2315: data = 9'o652;
		14'h2316: data = 9'o651;
		14'h2317: data = 9'o652;
		14'h2318: data = 9'o652;
		14'h2319: data = 9'o651;
		14'h231a: data = 9'o651;
		14'h231b: data = 9'o651;
		14'h231c: data = 9'o652;
		14'h231d: data = 9'o651;
		14'h231e: data = 9'o0;
		14'h231f: data = 9'o0;
		14'h2320: data = 9'o0;
		14'h2321: data = 9'o0;
		14'h2322: data = 9'o0;
		14'h2323: data = 9'o0;
		14'h2324: data = 9'o0;
		14'h2325: data = 9'o0;
		14'h2326: data = 9'o0;
		14'h2327: data = 9'o0;
		14'h2328: data = 9'o0;
		14'h2329: data = 9'o0;
		14'h232a: data = 9'o0;
		14'h232b: data = 9'o0;
		14'h232c: data = 9'o0;
		14'h232d: data = 9'o0;
		14'h232e: data = 9'o0;
		14'h232f: data = 9'o0;
		14'h2330: data = 9'o0;
		14'h2331: data = 9'o0;
		14'h2332: data = 9'o0;
		14'h2333: data = 9'o0;
		14'h2334: data = 9'o0;
		14'h2335: data = 9'o0;
		14'h2336: data = 9'o0;
		14'h2337: data = 9'o0;
		14'h2338: data = 9'o0;
		14'h2339: data = 9'o0;
		14'h233a: data = 9'o0;
		14'h233b: data = 9'o0;
		14'h233c: data = 9'o0;
		14'h233d: data = 9'o0;
		14'h233e: data = 9'o0;
		14'h233f: data = 9'o0;
		14'h2340: data = 9'o0;
		14'h2341: data = 9'o0;
		14'h2342: data = 9'o0;
		14'h2343: data = 9'o0;
		14'h2344: data = 9'o0;
		14'h2345: data = 9'o0;
		14'h2346: data = 9'o0;
		14'h2347: data = 9'o0;
		14'h2348: data = 9'o0;
		14'h2349: data = 9'o0;
		14'h234a: data = 9'o0;
		14'h234b: data = 9'o0;
		14'h234c: data = 9'o0;
		14'h234d: data = 9'o0;
		14'h234e: data = 9'o0;
		14'h234f: data = 9'o0;
		14'h2350: data = 9'o0;
		14'h2351: data = 9'o0;
		14'h2352: data = 9'o0;
		14'h2353: data = 9'o0;
		14'h2354: data = 9'o0;
		14'h2355: data = 9'o0;
		14'h2356: data = 9'o0;
		14'h2357: data = 9'o0;
		14'h2358: data = 9'o0;
		14'h2359: data = 9'o0;
		14'h235a: data = 9'o0;
		14'h235b: data = 9'o0;
		14'h235c: data = 9'o0;
		14'h235d: data = 9'o0;
		14'h235e: data = 9'o0;
		14'h235f: data = 9'o0;
		14'h2360: data = 9'o0;
		14'h2361: data = 9'o0;
		14'h2362: data = 9'o0;
		14'h2363: data = 9'o0;
		14'h2364: data = 9'o0;
		14'h2365: data = 9'o0;
		14'h2366: data = 9'o0;
		14'h2367: data = 9'o0;
		14'h2368: data = 9'o0;
		14'h2369: data = 9'o0;
		14'h236a: data = 9'o0;
		14'h236b: data = 9'o0;
		14'h236c: data = 9'o0;
		14'h236d: data = 9'o0;
		14'h236e: data = 9'o0;
		14'h236f: data = 9'o0;
		14'h2370: data = 9'o0;
		14'h2371: data = 9'o0;
		14'h2372: data = 9'o0;
		14'h2373: data = 9'o0;
		14'h2374: data = 9'o0;
		14'h2375: data = 9'o0;
		14'h2376: data = 9'o0;
		14'h2377: data = 9'o0;
		14'h2378: data = 9'o0;
		14'h2379: data = 9'o0;
		14'h237a: data = 9'o0;
		14'h237b: data = 9'o0;
		14'h237c: data = 9'o0;
		14'h237d: data = 9'o0;
		14'h237e: data = 9'o0;
		14'h237f: data = 9'o0;
		14'h2380: data = 9'o0;
		14'h2381: data = 9'o0;
		14'h2382: data = 9'o0;
		14'h2383: data = 9'o0;
		14'h2384: data = 9'o0;
		14'h2385: data = 9'o0;
		14'h2386: data = 9'o0;
		14'h2387: data = 9'o0;
		14'h2388: data = 9'o0;
		14'h2389: data = 9'o0;
		14'h238a: data = 9'o0;
		14'h238b: data = 9'o0;
		14'h238c: data = 9'o0;
		14'h238d: data = 9'o0;
		14'h238e: data = 9'o0;
		14'h238f: data = 9'o0;
		14'h2390: data = 9'o0;
		14'h2391: data = 9'o0;
		14'h2392: data = 9'o0;
		14'h2393: data = 9'o0;
		14'h2394: data = 9'o0;
		14'h2395: data = 9'o0;
		14'h2396: data = 9'o0;
		14'h2397: data = 9'o0;
		14'h2398: data = 9'o0;
		14'h2399: data = 9'o0;
		14'h239a: data = 9'o0;
		14'h239b: data = 9'o0;
		14'h239c: data = 9'o0;
		14'h239d: data = 9'o0;
		14'h239e: data = 9'o0;
		14'h239f: data = 9'o0;
		14'h23a0: data = 9'o0;
		14'h23a1: data = 9'o0;
		14'h23a2: data = 9'o0;
		14'h23a3: data = 9'o0;
		14'h23a4: data = 9'o0;
		14'h23a5: data = 9'o0;
		14'h23a6: data = 9'o0;
		14'h23a7: data = 9'o0;
		14'h23a8: data = 9'o0;
		14'h23a9: data = 9'o0;
		14'h23aa: data = 9'o0;
		14'h23ab: data = 9'o0;
		14'h23ac: data = 9'o0;
		14'h23ad: data = 9'o0;
		14'h23ae: data = 9'o0;
		14'h23af: data = 9'o0;
		14'h23b0: data = 9'o0;
		14'h23b1: data = 9'o0;
		14'h23b2: data = 9'o0;
		14'h23b3: data = 9'o0;
		14'h23b4: data = 9'o0;
		14'h23b5: data = 9'o0;
		14'h23b6: data = 9'o0;
		14'h23b7: data = 9'o0;
		14'h23b8: data = 9'o0;
		14'h23b9: data = 9'o0;
		14'h23ba: data = 9'o0;
		14'h23bb: data = 9'o0;
		14'h23bc: data = 9'o0;
		14'h23bd: data = 9'o0;
		14'h23be: data = 9'o0;
		14'h23bf: data = 9'o0;
		14'h23c0: data = 9'o0;
		14'h23c1: data = 9'o0;
		14'h23c2: data = 9'o0;
		14'h23c3: data = 9'o0;
		14'h23c4: data = 9'o0;
		14'h23c5: data = 9'o0;
		14'h23c6: data = 9'o0;
		14'h23c7: data = 9'o0;
		14'h23c8: data = 9'o0;
		14'h23c9: data = 9'o0;
		14'h23ca: data = 9'o0;
		14'h23cb: data = 9'o0;
		14'h23cc: data = 9'o0;
		14'h23cd: data = 9'o0;
		14'h23ce: data = 9'o0;
		14'h23cf: data = 9'o0;
		14'h23d0: data = 9'o0;
		14'h23d1: data = 9'o0;
		14'h23d2: data = 9'o0;
		14'h23d3: data = 9'o0;
		14'h23d4: data = 9'o0;
		14'h23d5: data = 9'o0;
		14'h23d6: data = 9'o0;
		14'h23d7: data = 9'o0;
		14'h23d8: data = 9'o0;
		14'h23d9: data = 9'o0;
		14'h23da: data = 9'o0;
		14'h23db: data = 9'o0;
		14'h23dc: data = 9'o0;
		14'h23dd: data = 9'o0;
		14'h23de: data = 9'o0;
		14'h23df: data = 9'o0;
		14'h23e0: data = 9'o0;
		14'h23e1: data = 9'o0;
		14'h23e2: data = 9'o0;
		14'h23e3: data = 9'o0;
		14'h23e4: data = 9'o0;
		14'h23e5: data = 9'o0;
		14'h23e6: data = 9'o0;
		14'h23e7: data = 9'o0;
		14'h23e8: data = 9'o0;
		14'h23e9: data = 9'o0;
		14'h23ea: data = 9'o0;
		14'h23eb: data = 9'o0;
		14'h23ec: data = 9'o0;
		14'h23ed: data = 9'o0;
		14'h23ee: data = 9'o0;
		14'h23ef: data = 9'o0;
		14'h23f0: data = 9'o0;
		14'h23f1: data = 9'o0;
		14'h23f2: data = 9'o0;
		14'h23f3: data = 9'o0;
		14'h23f4: data = 9'o0;
		14'h23f5: data = 9'o0;
		14'h23f6: data = 9'o0;
		14'h23f7: data = 9'o0;
		14'h23f8: data = 9'o0;
		14'h23f9: data = 9'o0;
		14'h23fa: data = 9'o0;
		14'h23fb: data = 9'o0;
		14'h23fc: data = 9'o0;
		14'h23fd: data = 9'o0;
		14'h23fe: data = 9'o0;
		14'h23ff: data = 9'o0;
		14'h2400: data = 9'o0;
		14'h2401: data = 9'o0;
		14'h2402: data = 9'o0;
		14'h2403: data = 9'o0;
		14'h2404: data = 9'o0;
		14'h2405: data = 9'o0;
		14'h2406: data = 9'o0;
		14'h2407: data = 9'o0;
		14'h2408: data = 9'o0;
		14'h2409: data = 9'o0;
		14'h240a: data = 9'o0;
		14'h240b: data = 9'o0;
		14'h240c: data = 9'o0;
		14'h240d: data = 9'o0;
		14'h240e: data = 9'o0;
		14'h240f: data = 9'o0;
		14'h2410: data = 9'o0;
		14'h2411: data = 9'o0;
		14'h2412: data = 9'o0;
		14'h2413: data = 9'o0;
		14'h2414: data = 9'o0;
		14'h2415: data = 9'o0;
		14'h2416: data = 9'o0;
		14'h2417: data = 9'o0;
		14'h2418: data = 9'o0;
		14'h2419: data = 9'o0;
		14'h241a: data = 9'o0;
		14'h241b: data = 9'o0;
		14'h241c: data = 9'o0;
		14'h241d: data = 9'o0;
		14'h241e: data = 9'o0;
		14'h241f: data = 9'o0;
		14'h2420: data = 9'o0;
		14'h2421: data = 9'o0;
		14'h2422: data = 9'o0;
		14'h2423: data = 9'o0;
		14'h2424: data = 9'o0;
		14'h2425: data = 9'o0;
		14'h2426: data = 9'o0;
		14'h2427: data = 9'o0;
		14'h2428: data = 9'o0;
		14'h2429: data = 9'o0;
		14'h242a: data = 9'o0;
		14'h242b: data = 9'o0;
		14'h242c: data = 9'o0;
		14'h242d: data = 9'o0;
		14'h242e: data = 9'o0;
		14'h242f: data = 9'o0;
		14'h2430: data = 9'o0;
		14'h2431: data = 9'o0;
		14'h2432: data = 9'o0;
		14'h2433: data = 9'o0;
		14'h2434: data = 9'o0;
		14'h2435: data = 9'o0;
		14'h2436: data = 9'o0;
		14'h2437: data = 9'o0;
		14'h2438: data = 9'o0;
		14'h2439: data = 9'o0;
		14'h243a: data = 9'o0;
		14'h243b: data = 9'o0;
		14'h243c: data = 9'o0;
		14'h243d: data = 9'o0;
		14'h243e: data = 9'o0;
		14'h243f: data = 9'o0;
		14'h2440: data = 9'o0;
		14'h2441: data = 9'o0;
		14'h2442: data = 9'o0;
		14'h2443: data = 9'o0;
		14'h2444: data = 9'o0;
		14'h2445: data = 9'o0;
		14'h2446: data = 9'o0;
		14'h2447: data = 9'o0;
		14'h2448: data = 9'o0;
		14'h2449: data = 9'o0;
		14'h244a: data = 9'o0;
		14'h244b: data = 9'o0;
		14'h244c: data = 9'o0;
		14'h244d: data = 9'o0;
		14'h244e: data = 9'o0;
		14'h244f: data = 9'o0;
		14'h2450: data = 9'o0;
		14'h2451: data = 9'o0;
		14'h2452: data = 9'o0;
		14'h2453: data = 9'o0;
		14'h2454: data = 9'o0;
		14'h2455: data = 9'o0;
		14'h2456: data = 9'o0;
		14'h2457: data = 9'o0;
		14'h2458: data = 9'o0;
		14'h2459: data = 9'o0;
		14'h245a: data = 9'o0;
		14'h245b: data = 9'o0;
		14'h245c: data = 9'o0;
		14'h245d: data = 9'o0;
		14'h245e: data = 9'o0;
		14'h245f: data = 9'o0;
		14'h2460: data = 9'o0;
		14'h2461: data = 9'o0;
		14'h2462: data = 9'o0;
		14'h2463: data = 9'o0;
		14'h2464: data = 9'o0;
		14'h2465: data = 9'o0;
		14'h2466: data = 9'o0;
		14'h2467: data = 9'o0;
		14'h2468: data = 9'o0;
		14'h2469: data = 9'o0;
		14'h246a: data = 9'o0;
		14'h246b: data = 9'o0;
		14'h246c: data = 9'o0;
		14'h246d: data = 9'o0;
		14'h246e: data = 9'o0;
		14'h246f: data = 9'o0;
		14'h2470: data = 9'o0;
		14'h2471: data = 9'o0;
		14'h2472: data = 9'o0;
		14'h2473: data = 9'o0;
		14'h2474: data = 9'o0;
		14'h2475: data = 9'o0;
		14'h2476: data = 9'o0;
		14'h2477: data = 9'o0;
		14'h2478: data = 9'o0;
		14'h2479: data = 9'o0;
		14'h247a: data = 9'o0;
		14'h247b: data = 9'o0;
		14'h247c: data = 9'o0;
		14'h247d: data = 9'o0;
		14'h247e: data = 9'o0;
		14'h247f: data = 9'o0;
		14'h2480: data = 9'o0;
		14'h2481: data = 9'o0;
		14'h2482: data = 9'o0;
		14'h2483: data = 9'o0;
		14'h2484: data = 9'o0;
		14'h2485: data = 9'o0;
		14'h2486: data = 9'o0;
		14'h2487: data = 9'o0;
		14'h2488: data = 9'o0;
		14'h2489: data = 9'o0;
		14'h248a: data = 9'o0;
		14'h248b: data = 9'o0;
		14'h248c: data = 9'o0;
		14'h248d: data = 9'o0;
		14'h248e: data = 9'o0;
		14'h248f: data = 9'o0;
		14'h2490: data = 9'o0;
		14'h2491: data = 9'o0;
		14'h2492: data = 9'o0;
		14'h2493: data = 9'o0;
		14'h2494: data = 9'o0;
		14'h2495: data = 9'o0;
		14'h2496: data = 9'o0;
		14'h2497: data = 9'o0;
		14'h2498: data = 9'o0;
		14'h2499: data = 9'o0;
		14'h249a: data = 9'o0;
		14'h249b: data = 9'o0;
		14'h249c: data = 9'o0;
		14'h249d: data = 9'o0;
		14'h249e: data = 9'o0;
		14'h249f: data = 9'o0;
		14'h24a0: data = 9'o0;
		14'h24a1: data = 9'o0;
		14'h24a2: data = 9'o0;
		14'h24a3: data = 9'o0;
		14'h24a4: data = 9'o0;
		14'h24a5: data = 9'o0;
		14'h24a6: data = 9'o0;
		14'h24a7: data = 9'o0;
		14'h24a8: data = 9'o0;
		14'h24a9: data = 9'o0;
		14'h24aa: data = 9'o0;
		14'h24ab: data = 9'o0;
		14'h24ac: data = 9'o0;
		14'h24ad: data = 9'o0;
		14'h24ae: data = 9'o0;
		14'h24af: data = 9'o0;
		14'h24b0: data = 9'o0;
		14'h24b1: data = 9'o0;
		14'h24b2: data = 9'o0;
		14'h24b3: data = 9'o0;
		14'h24b4: data = 9'o0;
		14'h24b5: data = 9'o0;
		14'h24b6: data = 9'o0;
		14'h24b7: data = 9'o0;
		14'h24b8: data = 9'o0;
		14'h24b9: data = 9'o0;
		14'h24ba: data = 9'o0;
		14'h24bb: data = 9'o0;
		14'h24bc: data = 9'o0;
		14'h24bd: data = 9'o0;
		14'h24be: data = 9'o0;
		14'h24bf: data = 9'o0;
		14'h24c0: data = 9'o0;
		14'h24c1: data = 9'o0;
		14'h24c2: data = 9'o0;
		14'h24c3: data = 9'o0;
		14'h24c4: data = 9'o0;
		14'h24c5: data = 9'o0;
		14'h24c6: data = 9'o0;
		14'h24c7: data = 9'o0;
		14'h24c8: data = 9'o0;
		14'h24c9: data = 9'o0;
		14'h24ca: data = 9'o0;
		14'h24cb: data = 9'o0;
		14'h24cc: data = 9'o0;
		14'h24cd: data = 9'o0;
		14'h24ce: data = 9'o0;
		14'h24cf: data = 9'o0;
		14'h24d0: data = 9'o0;
		14'h24d1: data = 9'o0;
		14'h24d2: data = 9'o0;
		14'h24d3: data = 9'o0;
		14'h24d4: data = 9'o0;
		14'h24d5: data = 9'o0;
		14'h24d6: data = 9'o0;
		14'h24d7: data = 9'o0;
		14'h24d8: data = 9'o0;
		14'h24d9: data = 9'o0;
		14'h24da: data = 9'o0;
		14'h24db: data = 9'o0;
		14'h24dc: data = 9'o0;
		14'h24dd: data = 9'o0;
		14'h24de: data = 9'o0;
		14'h24df: data = 9'o0;
		14'h24e0: data = 9'o0;
		14'h24e1: data = 9'o0;
		14'h24e2: data = 9'o0;
		14'h24e3: data = 9'o0;
		14'h24e4: data = 9'o0;
		14'h24e5: data = 9'o0;
		14'h24e6: data = 9'o0;
		14'h24e7: data = 9'o0;
		14'h24e8: data = 9'o0;
		14'h24e9: data = 9'o0;
		14'h24ea: data = 9'o0;
		14'h24eb: data = 9'o0;
		14'h24ec: data = 9'o0;
		14'h24ed: data = 9'o0;
		14'h24ee: data = 9'o0;
		14'h24ef: data = 9'o0;
		14'h24f0: data = 9'o0;
		14'h24f1: data = 9'o0;
		14'h24f2: data = 9'o0;
		14'h24f3: data = 9'o0;
		14'h24f4: data = 9'o0;
		14'h24f5: data = 9'o0;
		14'h24f6: data = 9'o0;
		14'h24f7: data = 9'o0;
		14'h24f8: data = 9'o0;
		14'h24f9: data = 9'o0;
		14'h24fa: data = 9'o0;
		14'h24fb: data = 9'o0;
		14'h24fc: data = 9'o0;
		14'h24fd: data = 9'o0;
		14'h24fe: data = 9'o0;
		14'h24ff: data = 9'o0;
		14'h2500: data = 9'o0;
		14'h2501: data = 9'o0;
		14'h2502: data = 9'o0;
		14'h2503: data = 9'o0;
		14'h2504: data = 9'o0;
		14'h2505: data = 9'o0;
		14'h2506: data = 9'o0;
		14'h2507: data = 9'o0;
		14'h2508: data = 9'o0;
		14'h2509: data = 9'o0;
		14'h250a: data = 9'o0;
		14'h250b: data = 9'o0;
		14'h250c: data = 9'o0;
		14'h250d: data = 9'o0;
		14'h250e: data = 9'o0;
		14'h250f: data = 9'o0;
		14'h2510: data = 9'o0;
		14'h2511: data = 9'o0;
		14'h2512: data = 9'o0;
		14'h2513: data = 9'o0;
		14'h2514: data = 9'o0;
		14'h2515: data = 9'o0;
		14'h2516: data = 9'o0;
		14'h2517: data = 9'o0;
		14'h2518: data = 9'o0;
		14'h2519: data = 9'o0;
		14'h251a: data = 9'o0;
		14'h251b: data = 9'o0;
		14'h251c: data = 9'o0;
		14'h251d: data = 9'o0;
		14'h251e: data = 9'o0;
		14'h251f: data = 9'o0;
		14'h2520: data = 9'o0;
		14'h2521: data = 9'o0;
		14'h2522: data = 9'o0;
		14'h2523: data = 9'o0;
		14'h2524: data = 9'o0;
		14'h2525: data = 9'o0;
		14'h2526: data = 9'o0;
		14'h2527: data = 9'o0;
		14'h2528: data = 9'o0;
		14'h2529: data = 9'o0;
		14'h252a: data = 9'o0;
		14'h252b: data = 9'o0;
		14'h252c: data = 9'o0;
		14'h252d: data = 9'o0;
		14'h252e: data = 9'o0;
		14'h252f: data = 9'o0;
		14'h2530: data = 9'o0;
		14'h2531: data = 9'o0;
		14'h2532: data = 9'o0;
		14'h2533: data = 9'o0;
		14'h2534: data = 9'o0;
		14'h2535: data = 9'o0;
		14'h2536: data = 9'o0;
		14'h2537: data = 9'o0;
		14'h2538: data = 9'o0;
		14'h2539: data = 9'o0;
		14'h253a: data = 9'o0;
		14'h253b: data = 9'o0;
		14'h253c: data = 9'o0;
		14'h253d: data = 9'o0;
		14'h253e: data = 9'o0;
		14'h253f: data = 9'o0;
		14'h2540: data = 9'o0;
		14'h2541: data = 9'o0;
		14'h2542: data = 9'o0;
		14'h2543: data = 9'o0;
		14'h2544: data = 9'o0;
		14'h2545: data = 9'o0;
		14'h2546: data = 9'o0;
		14'h2547: data = 9'o0;
		14'h2548: data = 9'o0;
		14'h2549: data = 9'o0;
		14'h254a: data = 9'o0;
		14'h254b: data = 9'o0;
		14'h254c: data = 9'o0;
		14'h254d: data = 9'o0;
		14'h254e: data = 9'o0;
		14'h254f: data = 9'o0;
		14'h2550: data = 9'o0;
		14'h2551: data = 9'o0;
		14'h2552: data = 9'o0;
		14'h2553: data = 9'o0;
		14'h2554: data = 9'o0;
		14'h2555: data = 9'o0;
		14'h2556: data = 9'o0;
		14'h2557: data = 9'o0;
		14'h2558: data = 9'o0;
		14'h2559: data = 9'o0;
		14'h255a: data = 9'o0;
		14'h255b: data = 9'o0;
		14'h255c: data = 9'o0;
		14'h255d: data = 9'o0;
		14'h255e: data = 9'o0;
		14'h255f: data = 9'o0;
		14'h2560: data = 9'o0;
		14'h2561: data = 9'o0;
		14'h2562: data = 9'o0;
		14'h2563: data = 9'o0;
		14'h2564: data = 9'o0;
		14'h2565: data = 9'o0;
		14'h2566: data = 9'o0;
		14'h2567: data = 9'o0;
		14'h2568: data = 9'o0;
		14'h2569: data = 9'o0;
		14'h256a: data = 9'o0;
		14'h256b: data = 9'o0;
		14'h256c: data = 9'o0;
		14'h256d: data = 9'o0;
		14'h256e: data = 9'o0;
		14'h256f: data = 9'o0;
		14'h2570: data = 9'o0;
		14'h2571: data = 9'o0;
		14'h2572: data = 9'o0;
		14'h2573: data = 9'o0;
		14'h2574: data = 9'o0;
		14'h2575: data = 9'o0;
		14'h2576: data = 9'o0;
		14'h2577: data = 9'o0;
		14'h2578: data = 9'o0;
		14'h2579: data = 9'o0;
		14'h257a: data = 9'o0;
		14'h257b: data = 9'o0;
		14'h257c: data = 9'o0;
		14'h257d: data = 9'o0;
		14'h257e: data = 9'o0;
		14'h257f: data = 9'o0;
		14'h2580: data = 9'o0;
		14'h2581: data = 9'o0;
		14'h2582: data = 9'o0;
		14'h2583: data = 9'o0;
		14'h2584: data = 9'o0;
		14'h2585: data = 9'o0;
		14'h2586: data = 9'o0;
		14'h2587: data = 9'o0;
		14'h2588: data = 9'o0;
		14'h2589: data = 9'o0;
		14'h258a: data = 9'o0;
		14'h258b: data = 9'o0;
		14'h258c: data = 9'o0;
		14'h258d: data = 9'o0;
		14'h258e: data = 9'o0;
		14'h258f: data = 9'o0;
		14'h2590: data = 9'o0;
		14'h2591: data = 9'o0;
		14'h2592: data = 9'o0;
		14'h2593: data = 9'o0;
		14'h2594: data = 9'o0;
		14'h2595: data = 9'o0;
		14'h2596: data = 9'o0;
		14'h2597: data = 9'o0;
		14'h2598: data = 9'o0;
		14'h2599: data = 9'o0;
		14'h259a: data = 9'o0;
		14'h259b: data = 9'o0;
		14'h259c: data = 9'o0;
		14'h259d: data = 9'o0;
		14'h259e: data = 9'o0;
		14'h259f: data = 9'o0;
		14'h25a0: data = 9'o0;
		14'h25a1: data = 9'o0;
		14'h25a2: data = 9'o0;
		14'h25a3: data = 9'o0;
		14'h25a4: data = 9'o0;
		14'h25a5: data = 9'o0;
		14'h25a6: data = 9'o0;
		14'h25a7: data = 9'o0;
		14'h25a8: data = 9'o0;
		14'h25a9: data = 9'o0;
		14'h25aa: data = 9'o0;
		14'h25ab: data = 9'o0;
		14'h25ac: data = 9'o0;
		14'h25ad: data = 9'o0;
		14'h25ae: data = 9'o0;
		14'h25af: data = 9'o0;
		14'h25b0: data = 9'o0;
		14'h25b1: data = 9'o0;
		14'h25b2: data = 9'o0;
		14'h25b3: data = 9'o0;
		14'h25b4: data = 9'o0;
		14'h25b5: data = 9'o0;
		14'h25b6: data = 9'o0;
		14'h25b7: data = 9'o0;
		14'h25b8: data = 9'o0;
		14'h25b9: data = 9'o0;
		14'h25ba: data = 9'o0;
		14'h25bb: data = 9'o0;
		14'h25bc: data = 9'o0;
		14'h25bd: data = 9'o0;
		14'h25be: data = 9'o0;
		14'h25bf: data = 9'o0;
		14'h25c0: data = 9'o0;
		14'h25c1: data = 9'o0;
		14'h25c2: data = 9'o0;
		14'h25c3: data = 9'o0;
		14'h25c4: data = 9'o0;
		14'h25c5: data = 9'o0;
		14'h25c6: data = 9'o0;
		14'h25c7: data = 9'o0;
		14'h25c8: data = 9'o0;
		14'h25c9: data = 9'o0;
		14'h25ca: data = 9'o0;
		14'h25cb: data = 9'o0;
		14'h25cc: data = 9'o0;
		14'h25cd: data = 9'o0;
		14'h25ce: data = 9'o0;
		14'h25cf: data = 9'o0;
		14'h25d0: data = 9'o0;
		14'h25d1: data = 9'o0;
		14'h25d2: data = 9'o0;
		14'h25d3: data = 9'o0;
		14'h25d4: data = 9'o0;
		14'h25d5: data = 9'o0;
		14'h25d6: data = 9'o0;
		14'h25d7: data = 9'o0;
		14'h25d8: data = 9'o0;
		14'h25d9: data = 9'o0;
		14'h25da: data = 9'o0;
		14'h25db: data = 9'o0;
		14'h25dc: data = 9'o0;
		14'h25dd: data = 9'o0;
		14'h25de: data = 9'o0;
		14'h25df: data = 9'o0;
		14'h25e0: data = 9'o0;
		14'h25e1: data = 9'o0;
		14'h25e2: data = 9'o0;
		14'h25e3: data = 9'o0;
		14'h25e4: data = 9'o0;
		14'h25e5: data = 9'o0;
		14'h25e6: data = 9'o0;
		14'h25e7: data = 9'o0;
		14'h25e8: data = 9'o0;
		14'h25e9: data = 9'o0;
		14'h25ea: data = 9'o0;
		14'h25eb: data = 9'o0;
		14'h25ec: data = 9'o0;
		14'h25ed: data = 9'o0;
		14'h25ee: data = 9'o0;
		14'h25ef: data = 9'o0;
		14'h25f0: data = 9'o0;
		14'h25f1: data = 9'o0;
		14'h25f2: data = 9'o0;
		14'h25f3: data = 9'o0;
		14'h25f4: data = 9'o0;
		14'h25f5: data = 9'o0;
		14'h25f6: data = 9'o0;
		14'h25f7: data = 9'o0;
		14'h25f8: data = 9'o0;
		14'h25f9: data = 9'o0;
		14'h25fa: data = 9'o0;
		14'h25fb: data = 9'o0;
		14'h25fc: data = 9'o0;
		14'h25fd: data = 9'o0;
		14'h25fe: data = 9'o0;
		14'h25ff: data = 9'o0;
		14'h2600: data = 9'o0;
		14'h2601: data = 9'o0;
		14'h2602: data = 9'o0;
		14'h2603: data = 9'o0;
		14'h2604: data = 9'o0;
		14'h2605: data = 9'o0;
		14'h2606: data = 9'o0;
		14'h2607: data = 9'o0;
		14'h2608: data = 9'o0;
		14'h2609: data = 9'o0;
		14'h260a: data = 9'o0;
		14'h260b: data = 9'o0;
		14'h260c: data = 9'o0;
		14'h260d: data = 9'o0;
		14'h260e: data = 9'o0;
		14'h260f: data = 9'o0;
		14'h2610: data = 9'o0;
		14'h2611: data = 9'o0;
		14'h2612: data = 9'o0;
		14'h2613: data = 9'o0;
		14'h2614: data = 9'o0;
		14'h2615: data = 9'o0;
		14'h2616: data = 9'o0;
		14'h2617: data = 9'o0;
		14'h2618: data = 9'o0;
		14'h2619: data = 9'o0;
		14'h261a: data = 9'o0;
		14'h261b: data = 9'o0;
		14'h261c: data = 9'o0;
		14'h261d: data = 9'o0;
		14'h261e: data = 9'o0;
		14'h261f: data = 9'o0;
		14'h2620: data = 9'o0;
		14'h2621: data = 9'o0;
		14'h2622: data = 9'o0;
		14'h2623: data = 9'o0;
		14'h2624: data = 9'o0;
		14'h2625: data = 9'o0;
		14'h2626: data = 9'o0;
		14'h2627: data = 9'o0;
		14'h2628: data = 9'o0;
		14'h2629: data = 9'o0;
		14'h262a: data = 9'o0;
		14'h262b: data = 9'o0;
		14'h262c: data = 9'o0;
		14'h262d: data = 9'o0;
		14'h262e: data = 9'o0;
		14'h262f: data = 9'o0;
		14'h2630: data = 9'o0;
		14'h2631: data = 9'o0;
		14'h2632: data = 9'o0;
		14'h2633: data = 9'o0;
		14'h2634: data = 9'o0;
		14'h2635: data = 9'o0;
		14'h2636: data = 9'o0;
		14'h2637: data = 9'o0;
		14'h2638: data = 9'o0;
		14'h2639: data = 9'o0;
		14'h263a: data = 9'o0;
		14'h263b: data = 9'o0;
		14'h263c: data = 9'o0;
		14'h263d: data = 9'o0;
		14'h263e: data = 9'o0;
		14'h263f: data = 9'o0;
		14'h2640: data = 9'o0;
		14'h2641: data = 9'o0;
		14'h2642: data = 9'o0;
		14'h2643: data = 9'o0;
		14'h2644: data = 9'o0;
		14'h2645: data = 9'o0;
		14'h2646: data = 9'o0;
		14'h2647: data = 9'o0;
		14'h2648: data = 9'o0;
		14'h2649: data = 9'o0;
		14'h264a: data = 9'o0;
		14'h264b: data = 9'o0;
		14'h264c: data = 9'o0;
		14'h264d: data = 9'o0;
		14'h264e: data = 9'o0;
		14'h264f: data = 9'o0;
		14'h2650: data = 9'o0;
		14'h2651: data = 9'o0;
		14'h2652: data = 9'o0;
		14'h2653: data = 9'o0;
		14'h2654: data = 9'o0;
		14'h2655: data = 9'o0;
		14'h2656: data = 9'o0;
		14'h2657: data = 9'o0;
		14'h2658: data = 9'o0;
		14'h2659: data = 9'o0;
		14'h265a: data = 9'o0;
		14'h265b: data = 9'o0;
		14'h265c: data = 9'o0;
		14'h265d: data = 9'o0;
		14'h265e: data = 9'o0;
		14'h265f: data = 9'o0;
		14'h2660: data = 9'o0;
		14'h2661: data = 9'o0;
		14'h2662: data = 9'o0;
		14'h2663: data = 9'o0;
		14'h2664: data = 9'o0;
		14'h2665: data = 9'o0;
		14'h2666: data = 9'o0;
		14'h2667: data = 9'o0;
		14'h2668: data = 9'o0;
		14'h2669: data = 9'o0;
		14'h266a: data = 9'o0;
		14'h266b: data = 9'o0;
		14'h266c: data = 9'o0;
		14'h266d: data = 9'o0;
		14'h266e: data = 9'o0;
		14'h266f: data = 9'o0;
		14'h2670: data = 9'o0;
		14'h2671: data = 9'o0;
		14'h2672: data = 9'o0;
		14'h2673: data = 9'o0;
		14'h2674: data = 9'o0;
		14'h2675: data = 9'o0;
		14'h2676: data = 9'o0;
		14'h2677: data = 9'o0;
		14'h2678: data = 9'o0;
		14'h2679: data = 9'o0;
		14'h267a: data = 9'o0;
		14'h267b: data = 9'o0;
		14'h267c: data = 9'o0;
		14'h267d: data = 9'o0;
		14'h267e: data = 9'o0;
		14'h267f: data = 9'o0;
		14'h2680: data = 9'o0;
		14'h2681: data = 9'o0;
		14'h2682: data = 9'o0;
		14'h2683: data = 9'o0;
		14'h2684: data = 9'o0;
		14'h2685: data = 9'o0;
		14'h2686: data = 9'o0;
		14'h2687: data = 9'o0;
		14'h2688: data = 9'o0;
		14'h2689: data = 9'o0;
		14'h268a: data = 9'o0;
		14'h268b: data = 9'o0;
		14'h268c: data = 9'o0;
		14'h268d: data = 9'o0;
		14'h268e: data = 9'o0;
		14'h268f: data = 9'o0;
		14'h2690: data = 9'o0;
		14'h2691: data = 9'o0;
		14'h2692: data = 9'o0;
		14'h2693: data = 9'o0;
		14'h2694: data = 9'o0;
		14'h2695: data = 9'o0;
		14'h2696: data = 9'o0;
		14'h2697: data = 9'o0;
		14'h2698: data = 9'o0;
		14'h2699: data = 9'o0;
		14'h269a: data = 9'o0;
		14'h269b: data = 9'o0;
		14'h269c: data = 9'o0;
		14'h269d: data = 9'o0;
		14'h269e: data = 9'o0;
		14'h269f: data = 9'o0;
		14'h26a0: data = 9'o0;
		14'h26a1: data = 9'o0;
		14'h26a2: data = 9'o0;
		14'h26a3: data = 9'o0;
		14'h26a4: data = 9'o0;
		14'h26a5: data = 9'o0;
		14'h26a6: data = 9'o0;
		14'h26a7: data = 9'o0;
		14'h26a8: data = 9'o0;
		14'h26a9: data = 9'o0;
		14'h26aa: data = 9'o0;
		14'h26ab: data = 9'o0;
		14'h26ac: data = 9'o0;
		14'h26ad: data = 9'o0;
		14'h26ae: data = 9'o0;
		14'h26af: data = 9'o0;
		14'h26b0: data = 9'o0;
		14'h26b1: data = 9'o0;
		14'h26b2: data = 9'o0;
		14'h26b3: data = 9'o0;
		14'h26b4: data = 9'o0;
		14'h26b5: data = 9'o0;
		14'h26b6: data = 9'o0;
		14'h26b7: data = 9'o0;
		14'h26b8: data = 9'o0;
		14'h26b9: data = 9'o0;
		14'h26ba: data = 9'o0;
		14'h26bb: data = 9'o0;
		14'h26bc: data = 9'o0;
		14'h26bd: data = 9'o0;
		14'h26be: data = 9'o0;
		14'h26bf: data = 9'o0;
		14'h26c0: data = 9'o0;
		14'h26c1: data = 9'o0;
		14'h26c2: data = 9'o0;
		14'h26c3: data = 9'o0;
		14'h26c4: data = 9'o0;
		14'h26c5: data = 9'o0;
		14'h26c6: data = 9'o0;
		14'h26c7: data = 9'o0;
		14'h26c8: data = 9'o0;
		14'h26c9: data = 9'o0;
		14'h26ca: data = 9'o0;
		14'h26cb: data = 9'o0;
		14'h26cc: data = 9'o0;
		14'h26cd: data = 9'o0;
		14'h26ce: data = 9'o0;
		14'h26cf: data = 9'o0;
		14'h26d0: data = 9'o0;
		14'h26d1: data = 9'o0;
		14'h26d2: data = 9'o0;
		14'h26d3: data = 9'o0;
		14'h26d4: data = 9'o0;
		14'h26d5: data = 9'o0;
		14'h26d6: data = 9'o0;
		14'h26d7: data = 9'o0;
		14'h26d8: data = 9'o0;
		14'h26d9: data = 9'o0;
		14'h26da: data = 9'o0;
		14'h26db: data = 9'o0;
		14'h26dc: data = 9'o0;
		14'h26dd: data = 9'o0;
		14'h26de: data = 9'o0;
		14'h26df: data = 9'o0;
		14'h26e0: data = 9'o0;
		14'h26e1: data = 9'o0;
		14'h26e2: data = 9'o0;
		14'h26e3: data = 9'o0;
		14'h26e4: data = 9'o0;
		14'h26e5: data = 9'o0;
		14'h26e6: data = 9'o0;
		14'h26e7: data = 9'o0;
		14'h26e8: data = 9'o0;
		14'h26e9: data = 9'o0;
		14'h26ea: data = 9'o0;
		14'h26eb: data = 9'o0;
		14'h26ec: data = 9'o0;
		14'h26ed: data = 9'o0;
		14'h26ee: data = 9'o0;
		14'h26ef: data = 9'o0;
		14'h26f0: data = 9'o0;
		14'h26f1: data = 9'o0;
		14'h26f2: data = 9'o0;
		14'h26f3: data = 9'o0;
		14'h26f4: data = 9'o0;
		14'h26f5: data = 9'o0;
		14'h26f6: data = 9'o0;
		14'h26f7: data = 9'o0;
		14'h26f8: data = 9'o0;
		14'h26f9: data = 9'o0;
		14'h26fa: data = 9'o0;
		14'h26fb: data = 9'o0;
		14'h26fc: data = 9'o0;
		14'h26fd: data = 9'o0;
		14'h26fe: data = 9'o0;
		14'h26ff: data = 9'o0;
		14'h2700: data = 9'o0;
		14'h2701: data = 9'o0;
		14'h2702: data = 9'o0;
		14'h2703: data = 9'o0;
		14'h2704: data = 9'o0;
		14'h2705: data = 9'o0;
		14'h2706: data = 9'o0;
		14'h2707: data = 9'o0;
		14'h2708: data = 9'o0;
		14'h2709: data = 9'o0;
		14'h270a: data = 9'o0;
		14'h270b: data = 9'o0;
		14'h270c: data = 9'o0;
		14'h270d: data = 9'o0;
		14'h270e: data = 9'o0;
		14'h270f: data = 9'o0;

		default: data = 9'o0;
	endcase
end

endmodule
