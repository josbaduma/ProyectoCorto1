`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:09:37 03/31/2016 
// Design Name: 
// Module Name:    ROM_TextBottom 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_TextBottom(
    input [7:0] addr,
    output reg [209:0] data
    );

always @* begin
	case(addr)
		8'h00: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h01: data = 200'b000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h02: data = 200'b000000000000000000000000000000000000011000000000000000000000011101111100000000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h03: data = 200'b000000000000000000000000000000000000011000000000000000000000011111000111000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h04: data = 200'b000000000000000000000000000000000000011000000000000000000000000000000011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h05: data = 200'b000000000000000000000000000000111110011001100011011111011111011000000001100000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h06: data = 200'b000000000000000000000000000001100111011001100011010011100111011000000001100000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h07: data = 200'b000000000000000000000000000001100011011001100011000001100011011000000001100000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h08: data = 200'b000000000000000000000000000001100011011001100011000001100011011000000001100000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h09: data = 200'b000000000000000000000000000001100011011001100011000001100011011000000011000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h0a: data = 200'b000000000000000000000000000001100111011001110110010011100011011011000111000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h0b: data = 200'b000000000000000000000000000000111110011001111110011111000011011001111110000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h0c: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h0d: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h0e: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;
		8'h0f: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h10: data = 200'b000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h11: data = 200'b000000000000000000000000000000000000000001100000000000000000000001111100000000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h12: data = 200'b000000000000000000000000000000000000000001100000000000000000000011000111000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h13: data = 200'b000000000000000000000000000000000000000001100000000000000000000000000011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h14: data = 200'b000000000000000000000000000001111101111101111110001111100110001100000001100000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h15: data = 200'b000000000000000000000000000011001110011101110111011000110110001100000001100000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h16: data = 200'b000000000000000000000000000011000110001101100011011000000110001100000001100000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h17: data = 200'b000000000000000000000000000011000110001101100011011111100110001100000001100000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h18: data = 200'b000000000000000000000000000011000110001101100011011000110110001100000011000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h19: data = 200'b000000000000000000000000000011001110001101110111011100110111011011000111000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h1a: data = 200'b000000000000000000000000000001111100001101111110011111100111111001111110000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h1b: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h1c: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h1d: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;
		8'h1e: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h1f: data = 200'b000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h20: data = 200'b000000000000000000000110000000000000000000000000000000000111000001111111110000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h21: data = 200'b000000000000000000000110000000000000000000000000000000000111000000001100000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h22: data = 200'b000000000000000000000110000000000000000000000000000000000000000000001100000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h23: data = 200'b000000000000001111100110011000110111111000111111001111100110111110001100000000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h24: data = 200'b000000000000011001110110011000110011011101100111011000110110001110001100000000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h25: data = 200'b000000000000011000110110011000110011001101100011011000000110000110001100000000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h26: data = 200'b000000000000011000110110011000110011011101100011011111100110000110001100000000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h27: data = 200'b000000000000011000110110011000110001111101100011011000110110000110001100000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h28: data = 200'b000000000000011001110110011101100000001101100011011100110110000110001100000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h29: data = 200'b000000000000001111100110011111100011111001100011011111100110000110001100000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h2a: data = 200'b000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h2b: data = 200'b000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h2c: data = 200'b000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;
		8'h2d: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h2e: data = 200'b000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h2f: data = 200'b000000000000000000000000000000000000000000001100000000000000000001111100000000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h30: data = 200'b000000000000000000000000000000000000000000001100000000000000000011000111000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h31: data = 200'b000000000000000000000000000000000000000000001100000000000000000110000011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h32: data = 200'b000000000000000000000000000000000000011111001100011111011000110110000001100000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h33: data = 200'b000000000000000000000000000000000000110011101100110001111100110110000001100000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h34: data = 200'b000000000000000000000000000000000000110001101100110000001101110110000001100000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h35: data = 200'b000000000000000000000000000000000000110001101100111111001101100110000001100000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h36: data = 200'b000000000000000000000000000000000000110001101100110001100111100110000011000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h37: data = 200'b000000000000000000000000000000000000110011101100111001100111000011000111000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h38: data = 200'b000000000000000000000000000000000000011111001100111111000111000001111110000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h39: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h3a: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h3b: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;
		8'h3c: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h3d: data = 200'b000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h3e: data = 200'b000000000110000000000000000000000000000000000000000000000000000000111111000000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h3f: data = 200'b000000000110000000000000000000000000000000000011000000000000000001110011000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h40: data = 200'b000000000110000000000000000000000000000000000011000000000000000001100011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h41: data = 200'b001111100110011000110111111000111111001111101111111111100011111001100011000000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h42: data = 200'b011001110110011000110011011101100111011000110011001001110110011100110011000000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h43: data = 200'b011000110110011000110011001101100011011000000011000000110110001100011111000000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h44: data = 200'b011000110110011000110011011101100011011111100011000000110111111100111011000000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h45: data = 200'b011000110110011000110001111101100011011000110011000000110000001100110011000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h46: data = 200'b011001110110011101100000001101100011011100110011001001110000011101100011000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h47: data = 200'b001111100110011111100011111001100011011111101111001111100111111001100011000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h48: data = 200'b000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h49: data = 200'b000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h4a: data = 200'b000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;
		8'h4b: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h4c: data = 200'b000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h4d: data = 200'b000000000000000000000000000000000000000000110000000000000000000000111111000000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h4e: data = 200'b000000000000000000000000000000000000000000110000000000000000000001110011000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h4f: data = 200'b000000000000000000000000000000000000000000110000000000000000000001100011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h50: data = 200'b000000000000000000000000000000111110001111110011111111110011111001100011000000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h51: data = 200'b000000000000000000000000000001100111011001110110011101110110011100110011000000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h52: data = 200'b000000000000000000000000000001100011011000110110011000110110001100011111000000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h53: data = 200'b000000000000000000000000000001100011011000110110011000110110001100111011000000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h54: data = 200'b000000000000000000000000000001100011011000110110011000110110001100110011000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h55: data = 200'b000000000000000000000000000001100111011001110110011000110110011101100011000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h56: data = 200'b000000000000000000000000000000111110001111110110011000110011111001100011000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h57: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h58: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h59: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;
		8'h5a: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h5b: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h5c: data = 200'b000000000000000000000000000000000000000000000000000000000000000011000011000000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h5d: data = 200'b000000000000000000000000000000000000000000000000000000000000000011000011000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h5e: data = 200'b000000000000000000000000000000000000000000000000000000000000000011000011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h5f: data = 200'b000000000011111000111111001111100111111000111110011001100111110011000011000000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h60: data = 200'b000000000110011101100111011001110011011101100011011011001100111011111111000000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h61: data = 200'b000000000110001101100011011000110011001101100000001111001100011011000011000000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h62: data = 200'b000000000110001101100011011000110011011101111110001110001111111011000011000000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h63: data = 200'b000000000110001101100011011000110001111101100011001111000000011011000011000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h64: data = 200'b000000000110011101100011011001110000001101110011011011100000111011000011000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h65: data = 200'b000000000011111001100011001111100011111001111110111001101111110011000011000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h66: data = 200'b000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h67: data = 200'b000000000000000000000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h68: data = 200'b000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;
		8'h69: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h6a: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h6b: data = 200'b000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h6c: data = 200'b000000000000000000000000000000000000000000000011000000000000000000110011000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h6d: data = 200'b000000000000000000000000000000000000000000000011000000000000000000110011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h6e: data = 200'b000000111110001111110011111001111110001111101111110111111001111100110011000000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h6f: data = 200'b000001100111011001110110011100110111011000110011001100111011001110110011000000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h70: data = 200'b000001100011011000110110001100110011011000000011001100011011000110011111000000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h71: data = 200'b000001100011011000110110001100110111011111100011001100011011111110000011000000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h72: data = 200'b000001100011011000110110001100011111011000110011001100011000000110000011000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h73: data = 200'b000001100111011000110110011100000011011100110011001100011000001110000011000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h74: data = 200'b000000111110011000110011111000111110011111101111001100011011111100000011000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h75: data = 200'b000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h76: data = 200'b000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h77: data = 200'b000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;
		8'h78: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h79: data = 200'b000000000000000000000000000000000110011000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000;
		8'h7a: data = 200'b000000000000000000000000000000000110011000000000000000000000000000111111000000000000000000110000000000000000000000000000001110000000000000000000000011000000000001111000000000000000000000000000000000001111111110;
		8'h7b: data = 200'b000000000000000000000000000000000110011000000000000000011000000000000011000000000000000000110000000000000000000000000000001110000000000000000000000011000000000011011100000000000000000000000000000000001110000110;
		8'h7c: data = 200'b000000000000000000000000000000000110011000000000000000011000000000000011000000000000000000110000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000110;
		8'h7d: data = 200'b000000000000000000000000001111100110011000111110111111111111111100000011000000110001111100111111000111110001111110011111001100111110011111000111110011000111110000011100000011111011111011000110111111001100000110;
		8'h7e: data = 200'b000000000000000000000000011000110110011001100111001110011000000110011111000000110011000110111011101100011011001110110011101100100111010011101100111011001100111001111000000110001100111011000110011011101100000110;
		8'h7f: data = 200'b000000000000000000000000011000000110011001100011000110011000001110000011000000000011000000110001101100000011000110110001101100000011000001101100011011001100011011100000000110000000011011000110011001101100111110;
		8'h80: data = 200'b000000000000000000000000011111100110011001111111000110011000111100000011000000000011111100110001101111110011000110110001101100000011000001101111111011001111111111000000000111111000011011000110011011101100000110;
		8'h81: data = 200'b000000000000000000000000011000110110011000000011000110011001100000000011000000000011000110110001101100011011000110110001101100000011000001100000011011000000011111000000000110001100011011000110001111101100000110;
		8'h82: data = 200'b000000000000000000000000011100110110011000000111000110011001100000000011000000110011100110111011101110011011000110110011101100100111010011100000111011000000111011001100000111001100011011101100000001101100000110;
		8'h83: data = 200'b000000000000000000000000011111100110011001111110000111111000111110111111000000110011111100111111001111110011000110011111001100111110011111001111110011001111110001111000000111111000011011111100011111001100000110;
		8'h84: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h85: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001100000000000;
		8'h86: data = 200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000;	
	endcase
end

endmodule
