`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:58:27 05/01/2016 
// Design Name: 
// Module Name:    ROM_CardC 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_CardC(
    input [6:0] addr,
    output reg [269:0] data
    );

always @* begin
	case(addr)
		7'h0: data = 270'b011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011;
		7'h1: data = 270'b011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011;
		7'h2: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h3: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h4: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h5: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h6: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h7: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h8: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h9: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'ha: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'hb: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'hc: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'hd: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'he: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'hf: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h10: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h11: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h12: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011111111111111111111111111111111011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h13: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011111111111111111111111111111111111111111111111011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h14: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h15: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h16: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h17: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h18: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h19: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h1a: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h1b: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h1c: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h1d: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h1e: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h1f: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h20: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h21: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h22: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h23: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h24: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111011011011011111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h25: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111011011011111111111111111111011011011111011011111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h26: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011011011011011111111111111111011111111111111011111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h27: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011011111111011011111111111011011111111111011011111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h28: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111011111111111011011111111111011111111111111011011111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h29: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111011111111111111011011111011011111111111011011111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h2a: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111011011111111111011011111011011111111111011011111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h2b: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111011011111111111011011011011111111111011011111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h2c: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111011011111111111011011011111111011011111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h2d: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111011011011111111011011011111011011111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h2e: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111011011011011011011011011011111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h2f: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011011011011011011111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h30: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111011011111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h31: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111011011111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h32: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111011011111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h33: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111011011111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h34: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011011111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h35: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011011111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h36: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111011111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h37: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h38: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h39: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h3a: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h3b: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h3c: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111011111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h3d: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111011111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h3e: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111011011011111111111111011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h3f: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h40: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h41: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h42: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h43: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h44: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h45: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h46: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h47: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011111111111111111111111011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h48: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h49: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h4a: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h4b: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h4c: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h4d: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h4e: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h4f: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h50: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h51: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h52: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h53: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h54: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h55: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h56: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h57: data = 270'b011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011;
		7'h58: data = 270'b011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011;
		7'h59: data = 270'b011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011;
		
		default: data = 270'b0;
	endcase
end
endmodule
