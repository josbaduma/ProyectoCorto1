`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:48:34 05/27/2016 
// Design Name: 
// Module Name:    ROM_Nave 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_Nave(
    input [5:0] addr,
    output reg [49:0] data
    );

always @* begin
	case(addr)
		6'h00: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h01: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h02: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h03: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h04: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h05: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h06: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h07: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h08: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h09: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h0a: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h0b: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h0c: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h0d: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h0e: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h0f: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h10: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h11: data = 50'b00000000000000000000000011000000000000000000000000;
		6'h12: data = 50'b00000000000000000000000111100000000000000000000000;
		6'h13: data = 50'b00000000000000000000000111100000000000000000000000;
		6'h14: data = 50'b00000000000000000000000111100000000000000000000000;
		6'h15: data = 50'b00000000000000000000000111100000000000000000000000;
		6'h16: data = 50'b00000000000111111111111111111111111111100000000000;
		6'h17: data = 50'b00000000000111111111111111111111111111100000000000;
		6'h18: data = 50'b00000000000111111111111111111111111111100000000000;
		6'h19: data = 50'b00000000000111111111111111111111111111100000000000;
		6'h1a: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h1b: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h1c: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h1d: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h1e: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h1f: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h20: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h21: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h22: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h23: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h24: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h25: data = 50'b00000001111111111111111111111111111111111110000000;
		6'h26: data = 50'b00000000000000000000000000000000000000000000000000;
		6'h27: data = 50'b00000000000000000000000000000000000000000000000000;
		
		default: data = 50'b0;
	endcase
end

endmodule
