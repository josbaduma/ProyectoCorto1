`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    06:44:38 05/09/2016 
// Design Name: 
// Module Name:    ROM_Text 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_Text(
    input [4:0] addr,
    output reg [107:0] data
    );

always @* begin
	case(addr)
		5'h0: data = 108'b000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000;
		5'h1: data = 108'b000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000;
		5'h2: data = 108'b000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000001111111111;
		5'h3: data = 108'b000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000001111111111;
		5'h4: data = 108'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001111;
		5'h5: data = 108'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001111;
		5'h6: data = 108'b111111111100000000111111110000000011111111000000001111111100000011110000111100000011111111000000111100001111;
		5'h7: data = 108'b111111111100000000111111110000000011111111000000001111111100000011110000111100000011111111000000111100001111;
		5'h8: data = 108'b000000001111000011110000000000000011110000000000111100001111000011111100111100001111000000000000111100001111;
		5'h9: data = 108'b000000001111000011110000000000000011110000000000111100001111000011111100111100001111000000000000111100001111;
		5'ha: data = 108'b000000001111000011110000000000000011110000000000111100001111000000000011111100001111000000000000001111111111;
		5'hb: data = 108'b000000001111000011110000000000000011110000000000111100001111000000000011111100001111000000000000001111111111;
		5'hc: data = 108'b001111111100000011111111110000000011110000000000111111111111000000000000111100001111111111000000000000001111;
		5'hd: data = 108'b001111111100000011111111110000000011110000000000111111111111000000000000111100001111111111000000000000001111;
		5'he: data = 108'b111100000000000011110000111100000011110000000000000000001111000000000000111100001111000011110000000000001111;
		5'hf: data = 108'b111100000000000011110000111100000011110000000000000000001111000000000000111100001111000011110000000000001111;
		5'h10: data = 108'b111100000000000011110000111100000011110000000000000000001111000000000000111100001111000011110000000000001111;
		5'h11: data = 108'b111100000000000011110000111100000011110000000000000000001111000000000000111100001111000011110000000000001111;
		5'h12: data = 108'b001111111111000011111111110000000011110000000000001111111100000000000000111100001111111111000000000000001111;
		5'h13: data = 108'b001111111111000011111111110000000011110000000000001111111100000000000000111100001111111111000000000000001111;
		5'h14: data = 108'b000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000;
		5'h15: data = 108'b000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000;
		5'h16: data = 108'b000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000;
		5'h17: data = 108'b000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000;
		5'h18: data = 108'b000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000;
		5'h19: data = 108'b000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000;
		
		default: data = 108'b0;
	endcase
end

endmodule
