`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:53:57 04/30/2016 
// Design Name: 
// Module Name:    ROM_CardA 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_CardA(
    input [6:0] addr,
    output reg [248:0] data
    );

always @* begin
	case(addr)
		7'h0: data = 249'b110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h1: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h2: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h3: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h4: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h5: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h6: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h7: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h8: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h9: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'ha: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'hb: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'hc: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100100100100100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'hd: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110110110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'he: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'hf: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111110100000100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h10: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h11: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111000100111111111111111111111111111111111000100100111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h12: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111100000100111111111111111111111111111111111100000100111111111111111111111111111111100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h13: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111100100000110111111111111111111111111111111000100000111111111111111111111111111111000100100110111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h14: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111110100100100100111111111111111111111111111111000000000111111111111111111111111111111000100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h15: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111100100100100100111111111111111111111111111111111111111111111111111111111111111111100000100100100110111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h16: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111100100100100100100111111111111111111111111111111111111111111111111111111111111111100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h17: data = 249'b111111111111111111111111111111111111111111111111111111111111111111100100100100100100100111111111111111100100100000100100000100100100100111111111111100100100000100100100111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h18: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100100100111111110100100100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h19: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100100111111111111110100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h1a: data = 249'b111111111111111111111111111111111111111111111111111111111111111111100100100100100100100000111111111110100100100111111111111111100100100111111111111100100100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h1b: data = 249'b111111111111111111111111111111111111111111111111111111111111111111100100100100100100100000111111111111100100100111111111111111100100100111111111111100100100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h1c: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100100100111111111111110100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h1d: data = 249'b110111111111111111111111111111111111111111111111111111111111111111110100100100100100100111111111111111100100100110111111111000100100100111111111111111100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h1e: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110100100100100100100111111111111111100000100100100100100100100100100111111111111111100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h1f: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110000110110110000100111111111111111111111111111111111111111111111111111111111111110000100111110100000111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h20: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111110111111111111100111100000000000100100100100100100100100100100100100000100111110100111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h21: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110111111111111111100111100000110111100100100100100100100100100100110110100100111111110111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h22: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110110111111111111100111100111111111111110100100100100100100000111111111111100111111100111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h23: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111000111111111100000111100111111111111111100100100100100100110111111111111100111111100111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h24: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111000100100100000100111100111111111111111100100100100100100100111111111111100111111100000100100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h25: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110100100100100100100111100100111111111100100100100100100100000111111111111100111110100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h26: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110100100100100100100111100100100100100100100100100100100100100100100100000100111110100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h27: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110100100100100100100111100100100000100100100100100100100100100100000100100100111110100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h28: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110100100100100100100111100100100100100100100100100100100100100100100100100100111110100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h29: data = 249'b111111111111111111111111111111111111111111111111111111111111111111110100100100100100100111100100100100100100100100100100100100100100100100100100111110100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h2a: data = 249'b110111111111111111111111111111111111111111111111111111111111111111110100100100100100100111100100100100100100100100100100100100100100100100100100111110100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h2b: data = 249'b110111111111111111111111111111111111111111111111111111111111111111111100100100100100100111100100100100100100100100100100100100100100100100100100111110100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h2c: data = 249'b110111111111111111111111111111111111111111111111111111111111111111111100100100100100100111100100100100100100100100100100100100100100100100100100111110100100100100100100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h2d: data = 249'b110111111111111111111111111111111111111000100111111111111110000111110100100100100100100111100100100100100100100100100100100100100100100100100100111110100100100100100100111110100111111111111111000111111111111111111111111111111111111111111111111111111;
		7'h2e: data = 249'b111111111111111111111111111111111111111100000111111111111100100111110100100100100100100111100100100100100100100100100100100100100100100100100100111111100100100100100100111100000111111111111111000111111111111111111111111111111111111111111111111111111;
		7'h2f: data = 249'b111111111111111111111111111111111111111000000111111111111100000111110100100100100100100111100000100100100100100100100100100100100100100100100100111110100100100100100100111100100111111111111111000111111111111111111111111111111111111111111111111111111;
		7'h30: data = 249'b111111111111111111111111111111111111111110111111111111111111110111111110110110110110110111111110110110110110110110110110110110110110110110110110111111110110110110110110111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		7'h31: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111110111111110111111111111111111111110111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h32: data = 249'b111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111110;
		7'h33: data = 249'b111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111110;
		7'h34: data = 249'b111111111111111111111111111111111111110100100100100100100100100100100100100100100100000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111110;
		7'h35: data = 249'b111111111111111111111111111111111111100100100100100100100100100100100100100100000110111110100100100100100100100100110111100100100100100100100000100111110100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111110;
		7'h36: data = 249'b111111111111111111111111111111111111100100100100100100100100100100100100100100100111111111111100100100100100100111111111111100100100100100100100111111111111100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111110;
		7'h37: data = 249'b111111111111111111111111111111111111100100100100100100100100100100100100100100111111111111111100100100100100100111111111111111100100100100100110111111111111100100100100100100100100100100100100100100110111111111111111111111111111111111111111111111110;
		7'h38: data = 249'b111111111111111111111111111111111111100100100100100100100100100100100100100100111111111111111100100100100100100111111111111111100100100100100111111111111111100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111110;
		7'h39: data = 249'b111111111111111111111111111111111111100100100100100100100100100100100100100100110111111111111000100100100100100111111111111110100100100100100110111111111111100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111110;
		7'h3a: data = 249'b111111111111111111111111111111111110100100100100100100100100100100100100100100100111111111110100100100100100100110111111111100100100100100100100111111111110100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111110;
		7'h3b: data = 249'b111111111111111111111111111111111110100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111110;
		7'h3c: data = 249'b111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111110;
		7'h3d: data = 249'b111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000100100100100100100100100100100100100100100100100100100100100100100100100100110111111111111111111111111111111111111111111110;
		7'h3e: data = 249'b111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111110;
		7'h3f: data = 249'b111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111110000100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111110;
		7'h40: data = 249'b111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111000100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111110;
		7'h41: data = 249'b111111111111111111111111111111110100100100100100100100100100100100100100100100100100100100100000110111111111111111111111111111111111111111100000100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111110;
		7'h42: data = 249'b111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111000100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111110;
		7'h43: data = 249'b111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111110100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111110;
		7'h44: data = 249'b111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100110111111111111111111111111111111111111111110;
		7'h45: data = 249'b111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100110111111111111111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111110;
		7'h46: data = 249'b111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111110;
		7'h47: data = 249'b111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111110;
		7'h48: data = 249'b111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111110;
		7'h49: data = 249'b111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100111111111111111111111111111111111111111110;
		7'h4a: data = 249'b111111111111111111111111111100100100100100100100100100100100100100100100100100100100100000111111111111111111111111111111111111111111111111111111100100100100100100100100100100100100100100100100100100100100100110111111111111111111111111111111111111110;
		7'h4b: data = 249'b111111111111111111111111111110110110100110110110110110110110110110110110110110110110110110111111111111111111111111111111111111111111111111111111111110110100100110110110110110110110110110110110110110110110110111111111111111111111111111111111111111111;
		7'h4c: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h4d: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h4e: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h4f: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h50: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h51: data = 249'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		7'h52: data = 249'b110110110110110110110110110110110110110111110111110111110110111110111110111110111111111111111111111111110111111111111111111111111111111110110110110110110110110110110110110110110110110110110110111111110110110111111110110111111111111111111111111110110;
		
		default: data = 249'b0;
	endcase
end

endmodule
