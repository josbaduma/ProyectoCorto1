`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:08:51 03/31/2016 
// Design Name: 
// Module Name:    ROM_TextTop 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_TextTop(
    input [7:0] addr,
    output reg [209:0] data
    );

always @* begin
	case(addr)
		8'h00: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h01: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h02: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h03: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h04: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000001110000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000;
		8'h05: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000001110011111111000000000000000001110000000000000000000000000000000001110000000000000000000000110000000000000111111000000000000000000000000;
		8'h06: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000001110000000000000000000000000000000001110000000000000000000000110000000000001110011100000000000000000000000;
		8'h07: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000001110000000000000000000000000000000001110000000000000000000000110000000000000000001110000000000000000000000;
		8'h08: data = 210'b000000000000000000000000000001111000001111100111111000110000110011111110000110000000111000000000111110001111111100000001111110000111110001111111011111100000111110000110000111110000000001110000000000000000000000;
		8'h09: data = 210'b000000000000000000000000000011001100011100110001111000110000110001110111000110000000111000000001100111001111001110000000011110001110011100001110011001110001100111000110001100111000000011100000000000000000000000;
		8'h0a: data = 210'b000000000000000000000000000000001110011000000000111000110000110001100011100110000000111000000011100011001110000110000000001110011100001100001110000000110011100011000110011100011000001111100000000000000000000000;
		8'h0b: data = 210'b000000000000000000000000000000001110111000000000011000110000110001100011100110011111111000000011000011101110000111000000000110011000001110001110000000111011000011100110011000011100111110000000000000000000000000;
		8'h0c: data = 210'b000000000000000000000000000000111100111000000000011000110000110001100011100110000000111000000011111111101110000111000000000110011000001110001110000000111011111111100110011111111101111000000000000000000000000000;
		8'h0d: data = 210'b000000000000000000000000000011110000111111100000011000110000110001110011000110000000111000000000000011101110000111000000000110011000001110001110000000111000000011100110000000011101110000000000000000000000000000;
		8'h0e: data = 210'b000000000000000000000000000011000000111000111000011000110000110000111111100110000000111000000000000011101110000111000000000110011000001110001110000000111000000011100110000000011101100000000000000000000000000000;
		8'h0f: data = 210'b000000000000000000000000000011000000111000111000011000111000110000000011100110000000111000000000000011101110000110000000000110011100001100001110000000110000000011100110000000011101110000000000000000000000000000;
		8'h10: data = 210'b000000000000000000000000000011100110111100111000011000111001110001111111100110000000111000000011000111001111001110000000000110001110011100001110011001110011000111000110011000111001110000110000000000000000000000;
		8'h11: data = 210'b000000000000000000000000000001111100111111110000011000111111100011100011000110000000111000000001111110001111111100000000000110000111111000111100011111100001111110000110001111110000011111100000000000000000000000;
		8'h12: data = 210'b000000000000000000000000000000000000000000000000000000000000000011000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h13: data = 210'b000000000000000000000000000000000000000000000000000000000000000011000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h14: data = 210'b000000000000000000000000000000000000000000000000000000000000000011100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h15: data = 210'b000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h16: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h17: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h18: data = 210'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase
end

endmodule
