`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:15:14 04/02/2016 
// Design Name: 
// Module Name:    ROM_TextFigure 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_TextFigure(
    input [8:0] addr,
    output reg [159:0] data
    );

always @* begin
	case(addr)
		9'h0: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h1: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h2: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000111100000000000000000000000;
		9'h3: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000111100000111111100000000000;
		9'h4: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000111100011111111110000000000;
		9'h5: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000111100001111100000000;
		9'h6: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000110000000111100000000;
		9'h7: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000011110000000;
		9'h8: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000111111100000001111000111100000011100000111111000001111101110000111100000000000001110000000;
		9'h9: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000011111111111000001111000111100000011100001111111110001111111110000111100000000000001111000000;
		9'ha: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000011110000111100001111000111100000011100011110001111000000111110000111100000000000001111000000;
		9'hb: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000111100000011100001111000111100000011100011000000111000000011110000111100000000000000111000000;
		9'hc: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000111000000011110001111000111100000011100000000000111100000001110000111100000000000000111000000;
		9'hd: data = 160'b0000000000000000000000000000000000000000000000000000000000000000001111000000001110001111000111100000011100000000000011100000001110000111100000000000000111000000;
		9'he: data = 160'b0000000000000000000000000000000000000000000000000000000000000000001111000000001110001111000111100000011100000000000011100000001110000111100000000000000111000000;
		9'hf: data = 160'b0000000000000000000000000000000000000000000000000000000000000000001111000000001110001111000111100000011100000000000011100000001110000111100000000000001111000000;
		9'h10: data = 160'b0000000000000000000000000000000000000000000000000000000000000000001111000000001110001111000111100000011100000000000011100000001110000111100000000000001111000000;
		9'h11: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000111000000001110001111000111100000011100000000000011100000001110000111100000000000001111000000;
		9'h12: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000111000000011110001111000111100000011100000000000111100000001110000111100000000000011110000000;
		9'h13: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000111100000011110001111000111110000111100011000000111100000001110000111100110000000011110000000;
		9'h14: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000011110000111100001111000111111000111100011110001111000000001110000111100111100001111100000000;
		9'h15: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000001111111111000001111000111111111111000001111111110000000001110000111100011111111111000000000;
		9'h16: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000011111100000001111000111101111110000000111111100000000001110000111100000111111100000000000;
		9'h17: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h18: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h19: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h1a: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h1b: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h1c: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h1d: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h1e: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h1f: data = 160'b0000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000;
		9'h20: data = 160'b0000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000;
		9'h21: data = 160'b0000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000111111100000000000;
		9'h22: data = 160'b0000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111100000000000000000000000000000000000000000000011111111110000000000;
		9'h23: data = 160'b0000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111100001111100000000;
		9'h24: data = 160'b0000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111100000000000000000000000000000000000000000000110000000111100000000;
		9'h25: data = 160'b0000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000011110000000;
		9'h26: data = 160'b0000000000000000000000000000000000111111100000001111011111100000000011111110001111101110000111101111110000000001111111000001111000000111000000000000001110000000;
		9'h27: data = 160'b0000000000000000000000000000000011111111111000001111111111110000001111111111101111111110000111111111111000000111111111110001111000000111000000000000001111000000;
		9'h28: data = 160'b0000000000000000000000000000000011110000111100001111110001111000001111000011100000111110000111111000111100000111100001110001111000000111000000000000001111000000;
		9'h29: data = 160'b0000000000000000000000000000000111100000011100001111100000111000011110000000000000011110000111110000011100001111000000000001111000000111000000000000000111000000;
		9'h2a: data = 160'b0000000000000000000000000000000111000000011110001111000000111100011110000000000000001110000111100000011110001111000000000001111000000111000000000000000111000000;
		9'h2b: data = 160'b0000000000000000000000000000001111000000001110001111000000011100011110000000000000001110000111100000001110001111000000000001111000000111000000000000000111000000;
		9'h2c: data = 160'b0000000000000000000000000000001111000000001110001111000000011100011111111100000000001110000111100000001110001111111110000001111000000111000000000000000111000000;
		9'h2d: data = 160'b0000000000000000000000000000001111000000001110001111000000011100011111111111000000001110000111100000001110001111111111100001111000000111000000000000001111000000;
		9'h2e: data = 160'b0000000000000000000000000000001111000000001110001111000000011100011110000111100000001110000111100000001110001111000011110001111000000111000000000000001111000000;
		9'h2f: data = 160'b0000000000000000000000000000000111000000001110001111000000011100011110000011100000001110000111100000001110001111000001110001111000000111000000000000001111000000;
		9'h30: data = 160'b0000000000000000000000000000000111000000011110001111000000111100011110000011100000001110000111100000011110001111000001110001111000000111000000000000011110000000;
		9'h31: data = 160'b0000000000000000000000000000000111100000011110001111100000111100011110000011100000001110000111110000011110001111000001110001111100001111000110000000011110000000;
		9'h32: data = 160'b0000000000000000000000000000000011110000111100001111110001111000011111000111100000001110000111111000111100001111100011110001111110001111000111100001111100000000;
		9'h33: data = 160'b0000000000000000000000000000000001111111111000001110111111110000011111111111000000001110000111011111111000001111111111100001111111111110000011111111111000000000;
		9'h34: data = 160'b0000000000000000000000000000000000011111100000001110011111100000011101111110000000001110000111001111110000001110111111000001111011111100000000111111100000000000;
		9'h35: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h36: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h37: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h38: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h39: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h3a: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h3b: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h3c: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h3d: data = 160'b0000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h3e: data = 160'b0000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000;
		9'h3f: data = 160'b0000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000001111000000000000111111111111111100000;
		9'h40: data = 160'b0000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000001111000000000000111111111111111100000;
		9'h41: data = 160'b0000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000;
		9'h42: data = 160'b0000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000;
		9'h43: data = 160'b0000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000;
		9'h44: data = 160'b0000000000000000000000000000000000000011111110000000111100011110000001110001111111111000000000111110011100000001111111000001111011111011100000000011100000000000;
		9'h45: data = 160'b0000000000000000000000000000000000001111111111100000111100011110000001110001111111111110000001111111111100000111111111110001111011111111100000000011100000000000;
		9'h46: data = 160'b0000000000000000000000000000000000001111000011110000111100011110000001110000011110001110000011110001111100000111100001110001111000001111100000000011100000000000;
		9'h47: data = 160'b0000000000000000000000000000000000011110000001110000111100011110000001110000011100001111000011100000111100001111000000000001111000000111100000000011100000000000;
		9'h48: data = 160'b0000000000000000000000000000000000011100000001111000111100011110000001110000111100000111000111100000011100001111000000000001111000000011100000000011100000000000;
		9'h49: data = 160'b0000000000000000000000000000000000111100000000111000111100011110000001110000111100000111000111100000011100001111000000000001111000000011100000000011100000000000;
		9'h4a: data = 160'b0000000000000000000000000000000000111100000000111000111100011110000001110000011100000111000111100000011100001111111110000001111000000011100000000011100000000000;
		9'h4b: data = 160'b0000000000000000000000000000000000111100000000111000111100011110000001110000011110001110000111100000011100001111111111100001111000000011100000000011100000000000;
		9'h4c: data = 160'b0000000000000000000000000000000000111100000000111000111100011110000001110000001111111110000111100000011100001111000011110001111000000011100000000011100000000000;
		9'h4d: data = 160'b0000000000000000000000000000000000011100000000111000111100011110000001110000000111111111000111100000011100001111000001110001111000000011100000000011100000000000;
		9'h4e: data = 160'b0000000000000000000000000000000000011100000001111000111100011110000001110000000000000111000111100000011100001111000001110001111000000011100000000011100000000000;
		9'h4f: data = 160'b0000000000000000000000000000000000011110000001111000111100011111000011110000000000000111000111100000011100001111000001110001111000000011100000000011100000000000;
		9'h50: data = 160'b0000000000000000000000000000000000001111000011110000111100011111100011110000001111111111000111100000011100001111100011110001111000000011100000000011100000000000;
		9'h51: data = 160'b0000000000000000000000000000000000000111111111100000111100011111111111100000111111111110000111100000011100001111111111100001111000000011100000000011100000000000;
		9'h52: data = 160'b0000000000000000000000000000000000000001111110000000111100011110111111000001111000001111000111100000011100001110111111000001111000000011100000000011100000000000;
		9'h53: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000001110000000111100000000000000000000000000000000000000000000000000000000000000000000000;
		9'h54: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000001110000000011100000000000000000000000000000000000000000000000000000000000000000000000;
		9'h55: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000001111000000111100000000000000000000000000000000000000000000000000000000000000000000000;
		9'h56: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100001111100000000000000000000000000000000000000000000000000000000000000000000000;
		9'h57: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h58: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h59: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h5a: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h5b: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h5c: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000;
		9'h5d: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000;
		9'h5e: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000001111111000000000000;
		9'h5f: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000111111111111000000000;
		9'h60: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000001111000001111100000000;
		9'h61: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000011110000000011110000000;
		9'h62: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000111100000000011110000000;
		9'h63: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000111100000011111110001110000000011100111100000000001111000000;
		9'h64: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000111100001111111111101111000000111100111000000000001111000000;
		9'h65: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000111100001111000011100111000000111100111000000000001111000000;
		9'h66: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001110000111100011110000000000111000000111001111000000000000111000000;
		9'h67: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000001111000111100011110000000000111100001111001111000000000000111000000;
		9'h68: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111000111100011110000000000011100001111001111000000000000111000000;
		9'h69: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111000111100011111111100000011110001110000111000000000000111000000;
		9'h6a: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111000111100011111111111000011110011110000111000000000001111000000;
		9'h6b: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111000111100011110000111100001110011100000111000000000001111000000;
		9'h6c: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111000111100011110000011100001111011100000111100000000001111000000;
		9'h6d: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000001111000111100011110000011100000111111100000011100000000011110000000;
		9'h6e: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001111000111100011110000011100000111111000000011110000000011110000000;
		9'h6f: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000011110000111100011111000111100000111111000000001111100001111100000000;
		9'h70: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000111100011111111111000000011111000000000111111111111000000000;
		9'h71: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000111100011101111110000000011110000000000001111111100000000000;
		9'h72: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h73: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h74: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h75: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h76: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h77: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h78: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h79: data = 160'b0000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h7a: data = 160'b0000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h7b: data = 160'b0000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000;
		9'h7c: data = 160'b0000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000111111111110000000;
		9'h7d: data = 160'b0000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000001111000001110000000;
		9'h7e: data = 160'b0000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000011110000001110000000;
		9'h7f: data = 160'b0000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000011110000001110000000;
		9'h80: data = 160'b0000000000000011111110000000111100011110000001110001111111111000000000111110011100000001111111000011111111110001111110000000000111111000000011110000001110000000;
		9'h81: data = 160'b0000000000001111111111100000111100011110000001110001111111111110000001111111111100000111111111110011111111110011111111100000011111111110000011110000001110000000;
		9'h82: data = 160'b0000000000001111000011110000111100011110000001110000011110001110000011110001111100000111100001110000001111000111100011110000111110001111000001110000001110000000;
		9'h83: data = 160'b0000000000011110000001110000111100011110000001110000011100001111000011100000111100001111000000000000001111000110000001110000111000000111000001111100001110000000;
		9'h84: data = 160'b0000000000011100000001111000111100011110000001110000111100000111000111100000011100001111000000000000001111000000000001111000111000000011100000111111111110000000;
		9'h85: data = 160'b0000000000111100000000111000111100011110000001110000111100000111000111100000011100001111000000000000001111000000000000111000111000000011100000001111111110000000;
		9'h86: data = 160'b0000000000111100000000111000111100011110000001110000011100000111000111100000011100001111111110000000001111000000000000111001111111111111100000111110001110000000;
		9'h87: data = 160'b0000000000111100000000111000111100011110000001110000011110001110000111100000011100001111111111100000001111000000000000111000111111111111100000111100001110000000;
		9'h88: data = 160'b0000000000111100000000111000111100011110000001110000001111111110000111100000011100001111000011110000001111000000000000111000000000000011100001111000001110000000;
		9'h89: data = 160'b0000000000011100000000111000111100011110000001110000000111111111000111100000011100001111000001110000001111000000000000111000000000000011100001111000001110000000;
		9'h8a: data = 160'b0000000000011100000001111000111100011110000001110000000000000111000111100000011100001111000001110000001111000000000001111000000000000111100011110000001110000000;
		9'h8b: data = 160'b0000000000011110000001111000111100011111000011110000000000000111000111100000011100001111000001110000001111000110000001111000000000000111100011110000001110000000;
		9'h8c: data = 160'b0000000000001111000011110000111100011111100011110000001111111111000111100000011100001111100011110000001110000111100011110000111000001111000011100000001110000000;
		9'h8d: data = 160'b0000000000000111111111100000111100011111111111100000111111111110000111100000011100001111111111100011111110000011111111100000111111111110000111100000001110000000;
		9'h8e: data = 160'b0000000000000001111110000000111100011110111111000001111000001111000111100000011100001110111111000011111100000001111111000000001111111000000111100000001110000000;
		9'h8f: data = 160'b0000000000000000000000000000000000000000000000000001110000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h90: data = 160'b0000000000000000000000000000000000000000000000000001110000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h91: data = 160'b0000000000000000000000000000000000000000000000000001111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h92: data = 160'b0000000000000000000000000000000000000000000000000000111100001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h93: data = 160'b0000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h94: data = 160'b0000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h95: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h96: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h97: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h98: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000;
		9'h99: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000;
		9'h9a: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000001111111110000000;
		9'h9b: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000111111111110000000;
		9'h9c: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000001111000001110000000;
		9'h9d: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000011110000001110000000;
		9'h9e: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000011110000001110000000;
		9'h9f: data = 160'b0000000000000000000000000000000000000000000000000000000000000000001111111000000000011111001110000000111110000111110011100000001111111000000011110000001110000000;
		9'ha0: data = 160'b0000000000000000000000000000000000000000000000000000000000000000111111111110000001111111111110000001111111101111111111100000111111111110000011110000001110000000;
		9'ha1: data = 160'b0000000000000000000000000000000000000000000000000000000000000000111100001111000001111001111110000011110011111110001111100000111100001111000001110000001110000000;
		9'ha2: data = 160'b0000000000000000000000000000000000000000000000000000000000000001111000000111000011110000011110000011100001111100000111100001111000000111000001111100001110000000;
		9'ha3: data = 160'b0000000000000000000000000000000000000000000000000000000000000001110000000111100011100000001110000111100000111100000011100001110000000111100000111111111110000000;
		9'ha4: data = 160'b0000000000000000000000000000000000000000000000000000000000000011110000000011100011100000001110000111100000011100000011100011110000000011100000001111111110000000;
		9'ha5: data = 160'b0000000000000000000000000000000000000000000000000000000000000011110000000011100111100000001110000111100000011100000011100011110000000011100000111110001110000000;
		9'ha6: data = 160'b0000000000000000000000000000000000000000000000000000000000000011110000000011100111100000001110000111100000011100000011100011110000000011100000111100001110000000;
		9'ha7: data = 160'b0000000000000000000000000000000000000000000000000000000000000011110000000011100111100000001110000111100000011100000011100011110000000011100001111000001110000000;
		9'ha8: data = 160'b0000000000000000000000000000000000000000000000000000000000000001110000000011100011100000001110000111100000011100000011100001110000000011100001111000001110000000;
		9'ha9: data = 160'b0000000000000000000000000000000000000000000000000000000000000001110000000111100011100000001110000111100000011100000011100001110000000111100011110000001110000000;
		9'haa: data = 160'b0000000000000000000000000000000000000000000000000000000000000001111000000111100011110000011110000111100000011100000011100001111000000111100011110000001110000000;
		9'hab: data = 160'b0000000000000000000000000000000000000000000000000000000000000000111100001111000001111000111110000111100000011100000011100000111100001111000011100000001110000000;
		9'hac: data = 160'b0000000000000000000000000000000000000000000000000000000000000000011111111110000000111111111110000111100000011100000011100000011111111110000111100000001110000000;
		9'had: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000111111000000000011111101110000111100000011100000011100000000111111000000111100000001110000000;
		9'hae: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'haf: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hb0: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hb1: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hb2: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hb3: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hb4: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hb5: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hb6: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001110000000;
		9'hb7: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001110000000;
		9'hb8: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001110000000;
		9'hb9: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001110000000;
		9'hba: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001110000000;
		9'hbb: data = 160'b0000000000000000000000000000011111110000000000111110011100000001111111000000111111111100000000011111110000111000000111100000111111000000001110000000001110000000;
		9'hbc: data = 160'b0000000000000000000000000001111111111100000001111111111100000111111111110000111111111111000001111111111100011100001111000011111111110000001110000000001110000000;
		9'hbd: data = 160'b0000000000000000000000000001111000011110000011110001111100000111100001111000001111000111000001111000011100011110001111000111110001111000001110000000001110000000;
		9'hbe: data = 160'b0000000000000000000000000011110000001110000011100000111100001111000000111000001110000111100011110000000000001110011110000111000000111000001110000000001110000000;
		9'hbf: data = 160'b0000000000000000000000000011100000001111000111100000011100001110000000111100011110000011100011110000000000001111011100000111000000011100001111111111111110000000;
		9'hc0: data = 160'b0000000000000000000000000111100000000111000111100000011100011110000000011100011110000011100011110000000000000111111100000111000000011100001111111111111110000000;
		9'hc1: data = 160'b0000000000000000000000000111100000000111000111100000011100011110000000011100001110000011100011111111100000000011111000001111111111111100001110000000001110000000;
		9'hc2: data = 160'b0000000000000000000000000111100000000111000111100000011100011110000000011100001111000111000011111111111000000011111000000111111111111100001110000000001110000000;
		9'hc3: data = 160'b0000000000000000000000000111100000000111000111100000011100011110000000011100000111111111000011110000111100000111111000000000000000011100001110000000001110000000;
		9'hc4: data = 160'b0000000000000000000000000011100000000111000111100000011100001110000000011100000011111111100011110000011100000111111100000000000000011100001110000000001110000000;
		9'hc5: data = 160'b0000000000000000000000000011100000001111000111100000011100001110000000111100000000000011100011110000011100001111011110000000000000111100001110000000001110000000;
		9'hc6: data = 160'b0000000000000000000000000011110000001111000111100000011100001111000000111100000000000011100011110000011100001110001110000000000000111100001110000000001110000000;
		9'hc7: data = 160'b0000000000000000000000000001111000011110000111100000011100000111100001111000000111111111100011111000111100011110001111000111000001111000001110000000001110000000;
		9'hc8: data = 160'b0000000000000000000000000000111111111100000111100000011100000011111111110000011111111111000011111111111000111100000111000111111111110000001110000000001110000000;
		9'hc9: data = 160'b0000000000000000000000000000001111110000000111100000011100000000111111000000111100000111100011101111110000111100000111100001111111000000001110000000001110000000;
		9'hca: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111000000011110000000000000000000000000000000000000000000000000000000000000000000000;
		9'hcb: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111000000001110000000000000000000000000000000000000000000000000000000000000000000000;
		9'hcc: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100000011110000000000000000000000000000000000000000000000000000000000000000000000;
		9'hcd: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000011110000111110000000000000000000000000000000000000000000000000000000000000000000000;
		9'hce: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000;
		9'hcf: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hd0: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hd1: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hd2: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hd3: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hd4: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hd5: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000;
		9'hd6: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111111111110000000;
		9'hd7: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000011111000011110000000;
		9'hd8: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000011110000011110000000;
		9'hd9: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000011100000011110000000;
		9'hda: data = 160'b0000000000000000001111111000000000011111001110000000111111100000011111111110000000001111111000011111111110000011111001110000000111111000000111100000011110000000;
		9'hdb: data = 160'b0000000000000000111111111110000000111111111110000011111111111000011111111111100000111111111110011111111110000111111111110000011111111110000111100000011110000000;
		9'hdc: data = 160'b0000000000000000111100001111000001111000111110000011110000111100000111100011100000111100001110000001111000001111000111110000111110001111000011100000011110000000;
		9'hdd: data = 160'b0000000000000001111000000111000001110000011110000111100000011100000111000011110001111000000000000001111000001110000011110000111000000111000011110000011110000000;
		9'hde: data = 160'b0000000000000001110000000111100011110000001110000111000000011110001111000001110001111000000000000001111000011110000001110000111000000011100001111000011110000000;
		9'hdf: data = 160'b0000000000000011110000000011100011110000001110001111000000001110001111000001110001111000000000000001111000011110000001110000111000000011100000111111111110000000;
		9'he0: data = 160'b0000000000000011110000000011100011110000001110001111000000001110000111000001110001111111110000000001111000011110000001110001111111111111100000001111111110000000;
		9'he1: data = 160'b0000000000000011110000000011100011110000001110001111000000001110000111100011100001111111111100000001111000011110000001110000111111111111100000000000011110000000;
		9'he2: data = 160'b0000000000000011110000000011100011110000001110001111000000001110000011111111100001111000011110000001111000011110000001110000000000000011100000000000011110000000;
		9'he3: data = 160'b0000000000000001110000000011100011110000001110000111000000001110000001111111110001111000001110000001111000011110000001110000000000000011100000000000011110000000;
		9'he4: data = 160'b0000000000000001110000000111100011110000001110000111000000011110000000000001110001111000001110000001111000011110000001110000000000000111100000000000011110000000;
		9'he5: data = 160'b0000000000000001111000000111100011110000001110000111100000011110000000000001110001111000001110000001111000011110000001110000000000000111100000000000011110000000;
		9'he6: data = 160'b0000000000000000111100001111000011110000001110000011110000111100000011111111110001111100011110000001110000011110000001110000111000001111000000000000011110000000;
		9'he7: data = 160'b0000000000000000011111111110000011110000001110000001111111111000001111111111100001111111111100011111110000011110000001110000111111111110000000000000011110000000;
		9'he8: data = 160'b0000000000000000000111111000000011110000001110000000011111100000011110000011110001110111111000011111100000011110000001110000001111111000000000000000011110000000;
		9'he9: data = 160'b0000000000000000000000000000000000000000000000000000000000000000011100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hea: data = 160'b0000000000000000000000000000000000000000000000000000000000000000011100000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'heb: data = 160'b0000000000000000000000000000000000000000000000000000000000000000011110000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hec: data = 160'b0000000000000000000000000000000000000000000000000000000000000000001111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hed: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hee: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hef: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hf0: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hf1: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hf2: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hf3: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000000000000000000000000000000000000000000000;
		9'hf4: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000000000000000000000000001111111111110000000;
		9'hf5: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000001111000000000000000001111111111110000000;
		9'hf6: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000001111000000000000000000000000011110000000;
		9'hf7: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000001111000000000000000000000000011110000000;
		9'hf8: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000111100011110000000000000000000000000000000001111000000000000000000000000011110000000;
		9'hf9: data = 160'b0000000000000000000000000000000000000000000000000000000000000000111111100000111100011110000001111110000011111011100011111111110001111111000000000000011110000000;
		9'hfa: data = 160'b0000000000000000000000000000000000000000000000000000000000000011111111111000111100011110000111111111100011111111100011111111110011111111100000000000011110000000;
		9'hfb: data = 160'b0000000000000000000000000000000000000000000000000000000000000011110000111000111100011110001111100011110000001111100000001111000011000011110000000000011110000000;
		9'hfc: data = 160'b0000000000000000000000000000000000000000000000000000000000000111100000000000111100011110001110000001110000000111100000001111000000000001110000000000011110000000;
		9'hfd: data = 160'b0000000000000000000000000000000000000000000000000000000000000111100000000000111100011110001110000000111000000011100000001111000000000001110000111111111110000000;
		9'hfe: data = 160'b0000000000000000000000000000000000000000000000000000000000000111100000000000111100011110001110000000111000000011100000001111000000000011110000111111111110000000;
		9'hff: data = 160'b0000000000000000000000000000000000000000000000000000000000000111111111000000111100011110011111111111111000000011100000001111000000011111100000000000011110000000;
		9'h100: data = 160'b0000000000000000000000000000000000000000000000000000000000000111111111110000111100011110001111111111111000000011100000001111000001111111000000000000011110000000;
		9'h101: data = 160'b0000000000000000000000000000000000000000000000000000000000000111100001111000111100011110000000000000111000000011100000001111000011111000000000000000011110000000;
		9'h102: data = 160'b0000000000000000000000000000000000000000000000000000000000000111100000111000111100011110000000000000111000000011100000001111000011100000000000000000011110000000;
		9'h103: data = 160'b0000000000000000000000000000000000000000000000000000000000000111100000111000111100011110000000000001111000000011100000001111000111100000000000000000011110000000;
		9'h104: data = 160'b0000000000000000000000000000000000000000000000000000000000000111100000111000111100011110000000000001111000000011100000001111000111100000000000000000011110000000;
		9'h105: data = 160'b0000000000000000000000000000000000000000000000000000000000000111110001111000111100011110001110000011110000000011100000001110000011110000110000000000011110000000;
		9'h106: data = 160'b0000000000000000000000000000000000000000000000000000000000000111111111110000111100011110001111111111100000000011100011111110000001111111110001111111111110000000;
		9'h107: data = 160'b0000000000000000000000000000000000000000000000000000000000000111011111100000111100011110000011111110000000000011100011111100000000111111100001111111111110000000;
		9'h108: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h109: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h10a: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h10b: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h10c: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		9'h10d: data = 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase
end

endmodule
