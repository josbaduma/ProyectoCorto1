`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:45:16 04/14/2016 
// Design Name: 
// Module Name:    DrawSystem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DrawSystem(
    input clk,
    input [9:0] HCount,
    input [9:0] VCount,
    output [2:0] rgb
    );


endmodule
