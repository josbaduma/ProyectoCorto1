`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:07:39 05/06/2016 
// Design Name: 
// Module Name:    ROM_Numero 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_Numero(
    input [7:0] addr,
    output reg [13:0] data
    );

always @* begin
	case(addr)
		8'h0: data = 14'b00000000000000;
		8'h1: data = 14'b00011111111000;
		8'h2: data = 14'b00011111111000;
		8'h3: data = 14'b01111000011110;
		8'h4: data = 14'b01111000011110;
		8'h5: data = 14'b01111110011110;
		8'h6: data = 14'b01111110011110;
		8'h7: data = 14'b01111110011110;
		8'h8: data = 14'b01111110011110;
		8'h9: data = 14'b01111000011110;
		8'ha: data = 14'b01111000011110;
		8'hb: data = 14'b01111001111110;
		8'hc: data = 14'b01111001111110;
		8'hd: data = 14'b01111001111110;
		8'he: data = 14'b01111001111110;
		8'hf: data = 14'b01111000011110;
		8'h10: data = 14'b01111000011110;
		8'h11: data = 14'b00011111111000;
		8'h12: data = 14'b00011111111000;
		8'h13: data = 14'b00000000000000;
		8'h14: data = 14'b00000000000000;
		8'h15: data = 14'b00011110000000;
		8'h16: data = 14'b00011110000000;
		8'h17: data = 14'b00011111100000;
		8'h18: data = 14'b00011111100000;
		8'h19: data = 14'b00011111111110;
		8'h1a: data = 14'b00011111111110;
		8'h1b: data = 14'b00011110000000;
		8'h1c: data = 14'b00011110000000;
		8'h1d: data = 14'b00011110000000;
		8'h1e: data = 14'b00011110000000;
		8'h1f: data = 14'b00011110000000;
		8'h20: data = 14'b00011110000000;
		8'h21: data = 14'b00011110000000;
		8'h22: data = 14'b00011110000000;
		8'h23: data = 14'b00011110000000;
		8'h24: data = 14'b00011110000000;
		8'h25: data = 14'b00011110000000;
		8'h26: data = 14'b00011110000000;
		8'h27: data = 14'b00000000000000;
		8'h28: data = 14'b00000000000000;
		8'h29: data = 14'b00011111111000;
		8'h2a: data = 14'b00011111111000;
		8'h2b: data = 14'b01111000011110;
		8'h2c: data = 14'b01111000011110;
		8'h2d: data = 14'b01111000011110;
		8'h2e: data = 14'b01111000011110;
		8'h2f: data = 14'b01111000000000;
		8'h30: data = 14'b01111000000000;
		8'h31: data = 14'b00011110000000;
		8'h32: data = 14'b00011110000000;
		8'h33: data = 14'b00000111100000;
		8'h34: data = 14'b00000111100000;
		8'h35: data = 14'b00000001111000;
		8'h36: data = 14'b00000001111000;
		8'h37: data = 14'b00000000011110;
		8'h38: data = 14'b00000000011110;
		8'h39: data = 14'b01111111111110;
		8'h3a: data = 14'b01111111111110;
		8'h3b: data = 14'b00000000000000;
		8'h3c: data = 14'b00000000000000;
		8'h3d: data = 14'b00011111111000;
		8'h3e: data = 14'b00011111111000;
		8'h3f: data = 14'b01111000011110;
		8'h40: data = 14'b01111000011110;
		8'h41: data = 14'b01111000011110;
		8'h42: data = 14'b01111000011110;
		8'h43: data = 14'b01111000000000;
		8'h44: data = 14'b01111000000000;
		8'h45: data = 14'b00011111100000;
		8'h46: data = 14'b00011111100000;
		8'h47: data = 14'b01111000000000;
		8'h48: data = 14'b01111000000000;
		8'h49: data = 14'b01111000011110;
		8'h4a: data = 14'b01111000011110;
		8'h4b: data = 14'b01111000011110;
		8'h4c: data = 14'b01111000011110;
		8'h4d: data = 14'b00011111111000;
		8'h4e: data = 14'b00011111111000;
		8'h4f: data = 14'b00000000000000;
		8'h50: data = 14'b00000000000000;
		8'h51: data = 14'b00000000111100;
		8'h52: data = 14'b00000000111100;
		8'h53: data = 14'b00000000111100;
		8'h54: data = 14'b00000000111100;
		8'h55: data = 14'b00111100111100;
		8'h56: data = 14'b00111100111100;
		8'h57: data = 14'b00111100111100;
		8'h58: data = 14'b00111100111100;
		8'h59: data = 14'b00111100111100;
		8'h5a: data = 14'b00111100111100;
		8'h5b: data = 14'b00111100001111;
		8'h5c: data = 14'b00111100001111;
		8'h5d: data = 14'b11111111111111;
		8'h5e: data = 14'b11111111111111;
		8'h5f: data = 14'b00111100000000;
		8'h60: data = 14'b00111100000000;
		8'h61: data = 14'b00111100000000;
		8'h62: data = 14'b00111100000000;
		8'h63: data = 14'b00000000000000;
		8'h64: data = 14'b00000000000000;
		8'h65: data = 14'b01111111111110;
		8'h66: data = 14'b01111111111110;
		8'h67: data = 14'b00000000011110;
		8'h68: data = 14'b00000000011110;
		8'h69: data = 14'b00000000011110;
		8'h6a: data = 14'b00000000011110;
		8'h6b: data = 14'b00000000011110;
		8'h6c: data = 14'b00000000011110;
		8'h6d: data = 14'b00011111111110;
		8'h6e: data = 14'b00011111111110;
		8'h6f: data = 14'b01111000000000;
		8'h70: data = 14'b01111000000000;
		8'h71: data = 14'b01111000000000;
		8'h72: data = 14'b01111000000000;
		8'h73: data = 14'b00011110000000;
		8'h74: data = 14'b00011110000000;
		8'h75: data = 14'b00000111111110;
		8'h76: data = 14'b00000111111110;
		8'h77: data = 14'b00000000000000;
		8'h78: data = 14'b00000000000000;
		8'h79: data = 14'b00011111100000;
		8'h7a: data = 14'b00011111100000;
		8'h7b: data = 14'b00000111100000;
		8'h7c: data = 14'b00000111100000;
		8'h7d: data = 14'b00000001111000;
		8'h7e: data = 14'b00000001111000;
		8'h7f: data = 14'b00011111111110;
		8'h80: data = 14'b00011111111110;
		8'h81: data = 14'b01111000011110;
		8'h82: data = 14'b01111000011110;
		8'h83: data = 14'b01111000011110;
		8'h84: data = 14'b01111000011110;
		8'h85: data = 14'b01111000011110;
		8'h86: data = 14'b01111000011110;
		8'h87: data = 14'b01111000011110;
		8'h88: data = 14'b01111000011110;
		8'h89: data = 14'b00011111111000;
		8'h8a: data = 14'b00011111111000;
		8'h8b: data = 14'b00000000000000;
		8'h8c: data = 14'b00000000000000;
		8'h8d: data = 14'b01111111111110;
		8'h8e: data = 14'b01111111111110;
		8'h8f: data = 14'b01111000000000;
		8'h90: data = 14'b01111000000000;
		8'h91: data = 14'b00011110000000;
		8'h92: data = 14'b00011110000000;
		8'h93: data = 14'b00011110000000;
		8'h94: data = 14'b00011110000000;
		8'h95: data = 14'b00000111100000;
		8'h96: data = 14'b00000111100000;
		8'h97: data = 14'b00000111100000;
		8'h98: data = 14'b00000111100000;
		8'h99: data = 14'b00000001111000;
		8'h9a: data = 14'b00000001111000;
		8'h9b: data = 14'b00000001111000;
		8'h9c: data = 14'b00000001111000;
		8'h9d: data = 14'b00000001111000;
		8'h9e: data = 14'b00000001111000;
		8'h9f: data = 14'b00000000000000;
		8'ha0: data = 14'b00000000000000;
		8'ha1: data = 14'b00011111111000;
		8'ha2: data = 14'b00011111111000;
		8'ha3: data = 14'b01111000011110;
		8'ha4: data = 14'b01111000011110;
		8'ha5: data = 14'b01111000011110;
		8'ha6: data = 14'b01111000011110;
		8'ha7: data = 14'b01111001111110;
		8'ha8: data = 14'b01111001111110;
		8'ha9: data = 14'b00011111111000;
		8'haa: data = 14'b00011111111000;
		8'hab: data = 14'b01111110011110;
		8'hac: data = 14'b01111110011110;
		8'had: data = 14'b01111000011110;
		8'hae: data = 14'b01111000011110;
		8'haf: data = 14'b01111000011110;
		8'hb0: data = 14'b01111000011110;
		8'hb1: data = 14'b00011111111000;
		8'hb2: data = 14'b00011111111000;
		8'hb3: data = 14'b00000000000000;
		
		default: data = 14'b00000000000000;
	endcase
end

endmodule
