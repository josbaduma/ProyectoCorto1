`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:25:47 03/30/2016 
// Design Name: 
// Module Name:    ROM_Text 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_Text(
    input [7:0] addr,
	 output reg [199:0] data
    );

always @* begin
	case(addr)
		8'h00: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h01: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h02: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h03: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h04: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h05: data = 200'b00000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000001110000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000;
		8'h06: data = 200'b00000000000000000011111100000000000001100000000000000000000001110000000000000000000000000000000001110000000000000000011111111001110000000000000000000000000000000000000000000000000000000000000000000000;
		8'h07: data = 200'b00000000000000000111001110000000000001100000000000000000000001110000000000000000000000000000000001110000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h08: data = 200'b00000000000000001110000000000000000001100000000000000000000001110000000000000000000000000000000001110000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h09: data = 200'b00000000000000001110000000001111100001100001111100000111111011111110001111100001111110000000111111110001111100000000011100000001100001111111001100001100011111100111110000011110000000000000000000000000;
		8'h0a: data = 200'b00000000000000000111000000011100110001100011100110001110011001110000111001110001111000000001110011110011100110000000011100000001100011101110001100001100011110001100111000110011000000000000000000000000;
		8'h0b: data = 200'b00000000000000000111110000011000111001100011000111001100000001110000110000111001110000000001100001110011000111000000011100000001100111000110001100001100011100000000011001110000000000000000000000000000;
		8'h0c: data = 200'b00000000000000000001111100111000011001100111000011011100000001110001110000011001100000000011100001110111000011000000011111111001100111000110001100001100011000000000011101110000000000000000000000000000;
		8'h0d: data = 200'b00000000000000000000011110111111111001100111111111011100000001110001110000011001100000000011100001110111111111000000011100000001100111000110001100001100011000000000011100111100000000000000000000000000;
		8'h0e: data = 200'b00000000000000000000001110111000000001100111000000011100000001110001110000011001100000000011100001110111000000000000011100000001100011001110001100001100011000000111111100001111000000000000000000000000;
		8'h0f: data = 200'b00000000000000000000000110111000000001100111000000011100000001110001110000011001100000000011100001110111000000000000011100000001100111111100001100001100011000011100011100000011000000000000000000000000;
		8'h10: data = 200'b00000000000000000000001110111000000001100111000000001100000001110000110000111001100000000001100001110111000000000000011100000001100111000000001100011100011000011100011100000011000000000000000000000000;
		8'h11: data = 200'b00000000000000001100001110011100011001100011100011001110011001110000111001110001100000000001110011110011100011000000011100000001100111111110001110011100011000011100111101100111000000000000000000000000;
		8'h12: data = 200'b00000000000000000111111000001111110001100001111110000111111000111100011111100001100000000000111111110001111110000000011100000001100011000111000111111100011000001111111100111110000000000000000000000000;
		8'h13: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011000000000000000000000000000000000000000000000000000000000000;
		8'h14: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011000000000000000000000000000000000000000000000000000000000000;
		8'h15: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111000000000000000000000000000000000000000000000000000000000000;
		8'h16: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000;
		8'h17: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'h18: data = 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase
end

endmodule
