`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:25:16 05/02/2016 
// Design Name: 
// Module Name:    ROM_Title 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ROM_Title(
    input [5:0] addr,
    output reg [215:0] data
    );

always @* begin
	case(addr)
		6'h0: data = 216'b111111110000000000001111111100001111111111111111111111110000000011111111000000000000111111110000000011111111111111110000000000001111111111111111111100000000000000001111111111111111000000000000000000001111111100000000;
		6'h1: data = 216'b111111110000000000001111111100001111111111111111111111110000000011111111000000000000111111110000000011111111111111110000000000001111111111111111111100000000000000001111111111111111000000000000000000001111111100000000;
		6'h2: data = 216'b111111110000000000001111111100001111111111111111111111110000000011111111000000000000111111110000000011111111111111110000000000001111111111111111111100000000000000001111111111111111000000000000000000001111111100000000;
		6'h3: data = 216'b111111110000000000001111111100001111111111111111111111110000000011111111000000000000111111110000000011111111111111110000000000001111111111111111111100000000000000001111111111111111000000000000000000001111111100000000;
		6'h4: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000000011111111111111110000;
		6'h5: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000000011111111111111110000;
		6'h6: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000000011111111111111110000;
		6'h7: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000000011111111111111110000;
		6'h8: data = 216'b111111111111000011111111111100001111111100000000000000000000000011111111111100001111111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h9: data = 216'b111111111111000011111111111100001111111100000000000000000000000011111111111100001111111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'ha: data = 216'b111111111111000011111111111100001111111100000000000000000000000011111111111100001111111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'hb: data = 216'b111111111111000011111111111100001111111100000000000000000000000011111111111100001111111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'hc: data = 216'b111111110000111100001111111100001111111100000000000000000000000011111111000011110000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'hd: data = 216'b111111110000111100001111111100001111111100000000000000000000000011111111000011110000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'he: data = 216'b111111110000111100001111111100001111111100000000000000000000000011111111000011110000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'hf: data = 216'b111111110000111100001111111100001111111100000000000000000000000011111111000011110000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h10: data = 216'b111111110000111100001111111100001111111111111111111100000000000011111111000011110000111111110000111111110000000011111111000000001111111111111111111100000000000000000000111111110000000000000000111111110000000011111111;
		6'h11: data = 216'b111111110000111100001111111100001111111111111111111100000000000011111111000011110000111111110000111111110000000011111111000000001111111111111111111100000000000000000000111111110000000000000000111111110000000011111111;
		6'h12: data = 216'b111111110000111100001111111100001111111111111111111100000000000011111111000011110000111111110000111111110000000011111111000000001111111111111111111100000000000000000000111111110000000000000000111111110000000011111111;
		6'h13: data = 216'b111111110000111100001111111100001111111111111111111100000000000011111111000011110000111111110000111111110000000011111111000000001111111111111111111100000000000000000000111111110000000000000000111111110000000011111111;
		6'h14: data = 216'b111111110000111100001111111100001111111100000000000000000000000011111111000011110000111111110000111111110000000011111111000000001111111100001111111100000000000000000000111111110000000000000000111111111111111111111111;
		6'h15: data = 216'b111111110000111100001111111100001111111100000000000000000000000011111111000011110000111111110000111111110000000011111111000000001111111100001111111100000000000000000000111111110000000000000000111111111111111111111111;
		6'h16: data = 216'b111111110000111100001111111100001111111100000000000000000000000011111111000011110000111111110000111111110000000011111111000000001111111100001111111100000000000000000000111111110000000000000000111111111111111111111111;
		6'h17: data = 216'b111111110000111100001111111100001111111100000000000000000000000011111111000011110000111111110000111111110000000011111111000000001111111100001111111100000000000000000000111111110000000000000000111111111111111111111111;
		6'h18: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h19: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h1a: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h1b: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h1c: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h1d: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h1e: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h1f: data = 216'b111111110000000000001111111100001111111100000000000000000000000011111111000000000000111111110000111111110000000011111111000000001111111100000000111111110000000000000000111111110000000000000000111111110000000011111111;
		6'h20: data = 216'b111111110000000000001111111100001111111111111111111111110000000011111111000000000000111111110000000011111111111111110000000000001111111100000000111111110000000000001111111111111111000000000000111111110000000011111111;
		6'h21: data = 216'b111111110000000000001111111100001111111111111111111111110000000011111111000000000000111111110000000011111111111111110000000000001111111100000000111111110000000000001111111111111111000000000000111111110000000011111111;
		6'h22: data = 216'b111111110000000000001111111100001111111111111111111111110000000011111111000000000000111111110000000011111111111111110000000000001111111100000000111111110000000000001111111111111111000000000000111111110000000011111111;
		6'h23: data = 216'b111111110000000000001111111100001111111111111111111111110000000011111111000000000000111111110000000011111111111111110000000000001111111100000000111111110000000000001111111111111111000000000000111111110000000011111111;
		
		default: data = 215'b0;
	endcase
end
endmodule
